module rv_regs(i_clk, i_reset_n, i_rs_valid, i_rs1, i_rs2, i_rd, i_write, i_data, o_data1, o_data2);
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0006_;
  wire _0008_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0135_;
  wire _0137_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire _1569_;
  wire _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire _1577_;
  wire _1578_;
  wire _1579_;
  wire _1580_;
  wire _1581_;
  wire _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire _1600_;
  wire _1601_;
  wire _1602_;
  wire _1603_;
  wire _1604_;
  wire _1605_;
  wire _1606_;
  wire _1607_;
  wire _1608_;
  wire _1609_;
  wire _1610_;
  wire _1611_;
  wire _1612_;
  wire _1613_;
  wire _1614_;
  wire _1615_;
  wire _1616_;
  wire _1617_;
  wire _1618_;
  wire _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire _1623_;
  wire _1624_;
  wire _1625_;
  wire _1626_;
  wire _1627_;
  wire _1628_;
  wire _1629_;
  wire _1630_;
  wire _1631_;
  wire _1632_;
  wire _1633_;
  wire _1634_;
  wire _1635_;
  wire _1636_;
  wire _1637_;
  wire _1638_;
  wire _1639_;
  wire _1640_;
  wire _1641_;
  wire _1642_;
  wire _1643_;
  wire _1644_;
  wire _1645_;
  wire _1646_;
  wire _1647_;
  wire _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire _1652_;
  wire _1653_;
  wire _1654_;
  wire _1655_;
  wire _1656_;
  wire _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire _1661_;
  wire _1662_;
  wire _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire _1673_;
  wire _1674_;
  wire _1675_;
  wire _1676_;
  wire _1677_;
  wire _1678_;
  wire _1679_;
  wire _1680_;
  wire _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire _1691_;
  wire _1692_;
  wire _1693_;
  wire _1694_;
  wire _1695_;
  wire _1696_;
  wire _1697_;
  wire _1698_;
  wire _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire _1710_;
  wire _1711_;
  wire _1712_;
  wire _1713_;
  wire _1714_;
  wire _1715_;
  wire _1716_;
  wire _1717_;
  wire _1718_;
  wire _1719_;
  wire _1720_;
  wire _1721_;
  wire _1722_;
  wire _1723_;
  wire _1724_;
  wire _1725_;
  wire _1726_;
  wire _1727_;
  wire _1728_;
  wire _1729_;
  wire _1730_;
  wire _1731_;
  wire _1732_;
  wire _1733_;
  wire _1734_;
  wire _1735_;
  wire _1736_;
  wire _1737_;
  wire _1738_;
  wire _1739_;
  wire _1740_;
  wire _1741_;
  wire _1742_;
  wire _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  wire _1750_;
  wire _1751_;
  wire _1752_;
  wire _1753_;
  wire _1754_;
  wire _1755_;
  wire _1756_;
  wire _1757_;
  wire _1758_;
  wire _1759_;
  wire _1760_;
  wire _1761_;
  wire _1762_;
  wire _1763_;
  wire _1764_;
  wire _1765_;
  wire _1766_;
  wire _1767_;
  wire _1768_;
  wire _1769_;
  wire _1770_;
  wire _1771_;
  wire _1772_;
  wire _1773_;
  wire _1774_;
  wire _1775_;
  wire _1776_;
  wire _1777_;
  wire _1778_;
  wire _1779_;
  wire _1780_;
  wire _1781_;
  wire _1782_;
  wire _1783_;
  wire _1784_;
  wire _1785_;
  wire _1786_;
  wire _1787_;
  wire _1788_;
  wire _1789_;
  wire _1790_;
  wire _1791_;
  wire _1792_;
  wire _1793_;
  wire _1794_;
  wire _1795_;
  wire _1796_;
  wire _1797_;
  wire _1798_;
  wire _1799_;
  wire _1800_;
  wire _1801_;
  wire _1802_;
  wire _1803_;
  wire _1804_;
  wire _1805_;
  wire _1806_;
  wire _1807_;
  wire _1808_;
  wire _1809_;
  wire _1810_;
  wire _1811_;
  wire _1812_;
  wire _1813_;
  wire _1814_;
  wire _1815_;
  wire _1816_;
  wire _1817_;
  wire _1818_;
  wire _1819_;
  wire _1820_;
  wire _1821_;
  wire _1822_;
  wire _1823_;
  wire _1824_;
  wire _1825_;
  wire _1826_;
  wire _1827_;
  wire _1828_;
  wire _1829_;
  wire _1830_;
  wire _1831_;
  wire _1832_;
  wire _1833_;
  wire _1834_;
  wire _1835_;
  wire _1836_;
  wire _1837_;
  wire _1838_;
  wire _1839_;
  wire _1840_;
  wire _1841_;
  wire _1842_;
  wire _1843_;
  wire _1844_;
  wire _1845_;
  wire _1846_;
  wire _1847_;
  wire _1848_;
  wire _1849_;
  wire _1850_;
  wire _1851_;
  wire _1852_;
  wire _1853_;
  wire _1854_;
  wire _1855_;
  wire _1856_;
  wire _1857_;
  wire _1858_;
  wire _1859_;
  wire _1860_;
  wire _1861_;
  wire _1862_;
  wire _1863_;
  wire _1864_;
  wire _1865_;
  wire _1866_;
  wire _1867_;
  wire _1868_;
  wire _1869_;
  wire _1870_;
  wire _1871_;
  wire _1872_;
  wire _1873_;
  wire _1874_;
  wire _1875_;
  wire _1876_;
  wire _1877_;
  wire _1878_;
  wire _1879_;
  wire _1880_;
  wire _1881_;
  wire _1882_;
  wire _1883_;
  wire _1884_;
  wire _1885_;
  wire _1886_;
  wire _1887_;
  wire _1888_;
  wire _1889_;
  wire _1890_;
  wire _1891_;
  wire _1892_;
  wire _1893_;
  wire _1894_;
  wire _1895_;
  wire _1896_;
  wire _1897_;
  wire _1898_;
  wire _1899_;
  wire _1900_;
  wire _1901_;
  wire _1902_;
  wire _1903_;
  wire _1904_;
  wire _1905_;
  wire _1906_;
  wire _1907_;
  wire _1908_;
  wire _1909_;
  wire _1910_;
  wire _1911_;
  wire _1912_;
  wire _1913_;
  wire _1914_;
  wire _1915_;
  wire _1916_;
  wire _1917_;
  wire _1918_;
  wire _1919_;
  wire _1920_;
  wire _1921_;
  wire _1922_;
  wire _1923_;
  wire _1924_;
  wire _1925_;
  wire _1926_;
  wire _1927_;
  wire _1928_;
  wire _1929_;
  wire _1930_;
  wire _1931_;
  wire _1932_;
  wire _1933_;
  wire _1934_;
  wire _1935_;
  wire _1936_;
  wire _1937_;
  wire _1938_;
  wire _1939_;
  wire _1940_;
  wire _1941_;
  wire _1942_;
  wire _1943_;
  wire _1944_;
  wire _1945_;
  wire _1946_;
  wire _1947_;
  wire _1948_;
  wire _1949_;
  wire _1950_;
  wire _1951_;
  wire _1952_;
  wire _1953_;
  wire _1954_;
  wire _1955_;
  wire _1956_;
  wire _1957_;
  wire _1958_;
  wire _1959_;
  wire _1960_;
  wire _1961_;
  wire _1962_;
  wire _1963_;
  wire _1964_;
  wire _1965_;
  wire _1966_;
  wire _1967_;
  wire _1968_;
  wire _1969_;
  wire _1970_;
  wire _1971_;
  wire _1972_;
  wire _1973_;
  wire _1974_;
  wire _1975_;
  wire _1976_;
  wire _1977_;
  wire _1978_;
  wire _1979_;
  wire _1980_;
  wire _1981_;
  wire _1982_;
  wire _1983_;
  wire _1984_;
  wire _1985_;
  wire _1986_;
  wire _1987_;
  wire _1988_;
  wire _1989_;
  wire _1990_;
  wire _1991_;
  wire _1992_;
  wire _1993_;
  wire _1994_;
  wire _1995_;
  wire _1996_;
  wire _1997_;
  wire _1998_;
  wire _1999_;
  wire _2000_;
  wire _2001_;
  wire _2002_;
  wire _2003_;
  wire _2004_;
  wire _2005_;
  wire _2006_;
  wire _2007_;
  wire _2008_;
  wire _2009_;
  wire _2010_;
  wire _2011_;
  wire _2012_;
  wire _2013_;
  wire _2014_;
  wire _2015_;
  wire _2016_;
  wire _2017_;
  wire _2018_;
  wire _2019_;
  wire _2020_;
  wire _2021_;
  wire _2022_;
  wire _2023_;
  wire _2024_;
  wire _2025_;
  wire _2026_;
  wire _2027_;
  wire _2028_;
  wire _2029_;
  wire _2030_;
  wire _2031_;
  wire _2032_;
  wire _2033_;
  wire _2034_;
  wire _2035_;
  wire _2036_;
  wire _2037_;
  wire _2038_;
  wire _2039_;
  wire _2040_;
  wire _2041_;
  wire _2042_;
  wire _2043_;
  wire _2044_;
  wire _2045_;
  wire _2046_;
  wire _2047_;
  wire _2048_;
  wire _2049_;
  wire _2050_;
  wire _2051_;
  wire _2052_;
  wire _2053_;
  wire _2054_;
  wire _2055_;
  wire _2056_;
  wire _2057_;
  wire _2058_;
  wire _2059_;
  wire _2060_;
  wire _2061_;
  wire _2062_;
  wire _2063_;
  wire _2064_;
  wire _2065_;
  wire _2066_;
  wire _2067_;
  wire _2068_;
  wire _2069_;
  wire _2070_;
  wire _2071_;
  wire _2072_;
  wire _2073_;
  wire _2074_;
  wire _2075_;
  wire _2076_;
  wire _2077_;
  wire _2078_;
  wire _2079_;
  wire _2080_;
  wire _2081_;
  wire _2082_;
  wire _2083_;
  wire _2084_;
  wire _2085_;
  wire _2086_;
  wire _2087_;
  wire _2088_;
  wire _2089_;
  wire _2090_;
  wire _2091_;
  wire _2092_;
  wire _2093_;
  wire _2094_;
  wire _2095_;
  wire _2096_;
  wire _2097_;
  wire _2098_;
  wire _2099_;
  wire _2100_;
  wire _2101_;
  wire _2102_;
  wire _2103_;
  wire _2104_;
  wire _2105_;
  wire _2106_;
  wire _2107_;
  wire _2108_;
  wire _2109_;
  wire _2110_;
  wire _2111_;
  wire _2112_;
  wire _2113_;
  wire _2114_;
  wire _2115_;
  wire _2116_;
  wire _2117_;
  wire _2118_;
  wire _2119_;
  wire _2120_;
  wire _2121_;
  wire _2122_;
  wire _2123_;
  wire _2124_;
  wire _2125_;
  wire _2126_;
  wire _2127_;
  wire _2128_;
  wire _2129_;
  wire _2130_;
  wire _2131_;
  wire _2132_;
  wire _2133_;
  wire _2134_;
  wire _2135_;
  wire _2136_;
  wire _2137_;
  wire _2138_;
  wire _2139_;
  wire _2140_;
  wire _2141_;
  wire _2142_;
  wire _2143_;
  wire _2144_;
  wire _2145_;
  wire _2146_;
  wire _2147_;
  wire _2148_;
  wire _2149_;
  wire _2150_;
  wire _2151_;
  wire _2152_;
  wire _2153_;
  wire _2154_;
  wire _2155_;
  wire _2156_;
  wire _2157_;
  wire _2158_;
  wire _2159_;
  wire _2160_;
  wire _2161_;
  wire _2162_;
  wire _2163_;
  wire _2164_;
  wire _2165_;
  wire _2166_;
  wire _2167_;
  wire _2168_;
  wire _2169_;
  wire _2170_;
  wire _2171_;
  wire _2172_;
  wire _2173_;
  wire _2174_;
  wire _2175_;
  wire _2176_;
  wire _2177_;
  wire _2178_;
  wire _2179_;
  wire _2180_;
  wire _2181_;
  wire _2182_;
  wire _2183_;
  wire _2184_;
  wire _2185_;
  wire _2186_;
  wire _2187_;
  wire _2188_;
  wire _2189_;
  wire _2190_;
  wire _2191_;
  wire _2192_;
  wire _2193_;
  wire _2194_;
  wire _2195_;
  wire _2196_;
  wire _2197_;
  wire _2198_;
  wire _2199_;
  wire _2200_;
  wire _2201_;
  wire _2202_;
  wire _2203_;
  wire _2204_;
  wire _2205_;
  wire _2206_;
  wire _2207_;
  wire _2208_;
  wire _2209_;
  wire _2210_;
  wire _2211_;
  wire _2212_;
  wire _2213_;
  wire _2214_;
  wire _2215_;
  wire _2216_;
  wire _2217_;
  wire _2218_;
  wire _2219_;
  wire _2220_;
  wire _2221_;
  wire _2222_;
  wire _2223_;
  wire _2224_;
  wire _2225_;
  wire _2226_;
  wire _2227_;
  wire _2228_;
  wire _2229_;
  wire _2230_;
  wire _2231_;
  wire _2232_;
  wire _2233_;
  wire _2234_;
  wire _2235_;
  wire _2236_;
  wire _2237_;
  wire _2238_;
  wire _2239_;
  wire _2240_;
  wire _2241_;
  wire _2242_;
  wire _2243_;
  wire _2244_;
  wire _2245_;
  wire _2246_;
  wire _2247_;
  wire _2248_;
  wire _2249_;
  wire _2250_;
  wire _2251_;
  wire _2252_;
  wire _2253_;
  wire _2254_;
  wire _2255_;
  wire _2256_;
  wire _2257_;
  wire _2258_;
  wire _2259_;
  wire _2260_;
  wire _2261_;
  wire _2262_;
  wire _2263_;
  wire _2264_;
  wire _2265_;
  wire _2266_;
  wire _2267_;
  wire _2268_;
  wire _2269_;
  wire _2270_;
  wire _2271_;
  wire _2272_;
  wire _2273_;
  wire _2274_;
  wire _2275_;
  wire _2276_;
  wire _2277_;
  wire _2278_;
  wire _2279_;
  wire _2280_;
  wire _2281_;
  wire _2282_;
  wire _2283_;
  wire w_wr_sel_rd4;
  wire w_wr_sel_nrd4;
  wire _2285_;
  wire _2286_;
  wire _2287_;
  wire _2288_;
  wire _2289_;
  wire _2290_;
  wire _2291_;
  wire _2293_;
  wire _2294_;
  wire _2295_;
  wire _2296_;
  wire _2297_;
  wire w_wr_sel_nrd4_rd0_or_rd1;
  wire w_wr_sel_rd4_rd0_or_rd1;
  wire \g_bit[0].g_word[10].r_bit.DE ;
  wire \g_bit[0].g_word[10].r_bit.Q ;
  wire \g_bit[0].g_word[11].r_bit.DE ;
  wire \g_bit[0].g_word[11].r_bit.Q ;
  wire \g_bit[0].g_word[12].r_bit.DE ;
  wire \g_bit[0].g_word[12].r_bit.Q ;
  wire \g_bit[0].g_word[13].r_bit.DE ;
  wire \g_bit[0].g_word[13].r_bit.Q ;
  wire \g_bit[0].g_word[14].r_bit.DE ;
  wire \g_bit[0].g_word[14].r_bit.Q ;
  wire \g_bit[0].g_word[15].r_bit.DE ;
  wire \g_bit[0].g_word[15].r_bit.Q ;
  wire \g_bit[0].g_word[16].r_bit.DE ;
  wire \g_bit[0].g_word[16].r_bit.Q ;
  wire \g_bit[0].g_word[17].r_bit.DE ;
  wire \g_bit[0].g_word[17].r_bit.Q ;
  wire \g_bit[0].g_word[18].r_bit.DE ;
  wire \g_bit[0].g_word[18].r_bit.Q ;
  wire \g_bit[0].g_word[19].r_bit.DE ;
  wire \g_bit[0].g_word[19].r_bit.Q ;
  wire \g_bit[0].g_word[1].r_bit.DE ;
  wire \g_bit[0].g_word[1].r_bit.Q ;
  wire \g_bit[0].g_word[20].r_bit.DE ;
  wire \g_bit[0].g_word[20].r_bit.Q ;
  wire \g_bit[0].g_word[21].r_bit.DE ;
  wire \g_bit[0].g_word[21].r_bit.Q ;
  wire \g_bit[0].g_word[22].r_bit.DE ;
  wire \g_bit[0].g_word[22].r_bit.Q ;
  wire \g_bit[0].g_word[23].r_bit.DE ;
  wire \g_bit[0].g_word[23].r_bit.Q ;
  wire \g_bit[0].g_word[24].r_bit.DE ;
  wire \g_bit[0].g_word[24].r_bit.Q ;
  wire \g_bit[0].g_word[25].r_bit.DE ;
  wire \g_bit[0].g_word[25].r_bit.Q ;
  wire \g_bit[0].g_word[26].r_bit.DE ;
  wire \g_bit[0].g_word[26].r_bit.Q ;
  wire \g_bit[0].g_word[27].r_bit.DE ;
  wire \g_bit[0].g_word[27].r_bit.Q ;
  wire \g_bit[0].g_word[28].r_bit.DE ;
  wire \g_bit[0].g_word[28].r_bit.Q ;
  wire \g_bit[0].g_word[29].r_bit.DE ;
  wire \g_bit[0].g_word[29].r_bit.Q ;
  wire \g_bit[0].g_word[2].r_bit.DE ;
  wire \g_bit[0].g_word[2].r_bit.Q ;
  wire \g_bit[0].g_word[30].r_bit.DE ;
  wire \g_bit[0].g_word[30].r_bit.Q ;
  wire \g_bit[0].g_word[31].r_bit.DE ;
  wire \g_bit[0].g_word[31].r_bit.Q ;
  wire \g_bit[0].g_word[3].r_bit.DE ;
  wire \g_bit[0].g_word[3].r_bit.Q ;
  wire \g_bit[0].g_word[4].r_bit.DE ;
  wire \g_bit[0].g_word[4].r_bit.Q ;
  wire \g_bit[0].g_word[5].r_bit.DE ;
  wire \g_bit[0].g_word[5].r_bit.Q ;
  wire \g_bit[0].g_word[6].r_bit.DE ;
  wire \g_bit[0].g_word[6].r_bit.Q ;
  wire \g_bit[0].g_word[7].r_bit.DE ;
  wire \g_bit[0].g_word[7].r_bit.Q ;
  wire \g_bit[0].g_word[8].r_bit.DE ;
  wire \g_bit[0].g_word[8].r_bit.Q ;
  wire \g_bit[0].g_word[9].r_bit.DE ;
  wire \g_bit[0].g_word[9].r_bit.Q ;
  wire \g_bit[0].r_rs1.D ;
  wire \g_bit[0].r_rs1.Q ;
  wire \g_bit[0].r_rs2.D ;
  wire \g_bit[0].r_rs2.Q ;
  wire \g_bit[10].g_word[10].r_bit.Q ;
  wire \g_bit[10].g_word[11].r_bit.Q ;
  wire \g_bit[10].g_word[12].r_bit.Q ;
  wire \g_bit[10].g_word[13].r_bit.Q ;
  wire \g_bit[10].g_word[14].r_bit.Q ;
  wire \g_bit[10].g_word[15].r_bit.Q ;
  wire \g_bit[10].g_word[16].r_bit.Q ;
  wire \g_bit[10].g_word[17].r_bit.Q ;
  wire \g_bit[10].g_word[18].r_bit.Q ;
  wire \g_bit[10].g_word[19].r_bit.Q ;
  wire \g_bit[10].g_word[1].r_bit.Q ;
  wire \g_bit[10].g_word[20].r_bit.Q ;
  wire \g_bit[10].g_word[21].r_bit.Q ;
  wire \g_bit[10].g_word[22].r_bit.Q ;
  wire \g_bit[10].g_word[23].r_bit.Q ;
  wire \g_bit[10].g_word[24].r_bit.Q ;
  wire \g_bit[10].g_word[25].r_bit.Q ;
  wire \g_bit[10].g_word[26].r_bit.Q ;
  wire \g_bit[10].g_word[27].r_bit.Q ;
  wire \g_bit[10].g_word[28].r_bit.Q ;
  wire \g_bit[10].g_word[29].r_bit.Q ;
  wire \g_bit[10].g_word[2].r_bit.Q ;
  wire \g_bit[10].g_word[30].r_bit.Q ;
  wire \g_bit[10].g_word[31].r_bit.Q ;
  wire \g_bit[10].g_word[3].r_bit.Q ;
  wire \g_bit[10].g_word[4].r_bit.Q ;
  wire \g_bit[10].g_word[5].r_bit.Q ;
  wire \g_bit[10].g_word[6].r_bit.Q ;
  wire \g_bit[10].g_word[7].r_bit.Q ;
  wire \g_bit[10].g_word[8].r_bit.Q ;
  wire \g_bit[10].g_word[9].r_bit.Q ;
  wire \g_bit[10].r_rs1.D ;
  wire \g_bit[10].r_rs1.Q ;
  wire \g_bit[10].r_rs2.D ;
  wire \g_bit[10].r_rs2.Q ;
  wire \g_bit[11].g_word[10].r_bit.Q ;
  wire \g_bit[11].g_word[11].r_bit.Q ;
  wire \g_bit[11].g_word[12].r_bit.Q ;
  wire \g_bit[11].g_word[13].r_bit.Q ;
  wire \g_bit[11].g_word[14].r_bit.Q ;
  wire \g_bit[11].g_word[15].r_bit.Q ;
  wire \g_bit[11].g_word[16].r_bit.Q ;
  wire \g_bit[11].g_word[17].r_bit.Q ;
  wire \g_bit[11].g_word[18].r_bit.Q ;
  wire \g_bit[11].g_word[19].r_bit.Q ;
  wire \g_bit[11].g_word[1].r_bit.Q ;
  wire \g_bit[11].g_word[20].r_bit.Q ;
  wire \g_bit[11].g_word[21].r_bit.Q ;
  wire \g_bit[11].g_word[22].r_bit.Q ;
  wire \g_bit[11].g_word[23].r_bit.Q ;
  wire \g_bit[11].g_word[24].r_bit.Q ;
  wire \g_bit[11].g_word[25].r_bit.Q ;
  wire \g_bit[11].g_word[26].r_bit.Q ;
  wire \g_bit[11].g_word[27].r_bit.Q ;
  wire \g_bit[11].g_word[28].r_bit.Q ;
  wire \g_bit[11].g_word[29].r_bit.Q ;
  wire \g_bit[11].g_word[2].r_bit.Q ;
  wire \g_bit[11].g_word[30].r_bit.Q ;
  wire \g_bit[11].g_word[31].r_bit.Q ;
  wire \g_bit[11].g_word[3].r_bit.Q ;
  wire \g_bit[11].g_word[4].r_bit.Q ;
  wire \g_bit[11].g_word[5].r_bit.Q ;
  wire \g_bit[11].g_word[6].r_bit.Q ;
  wire \g_bit[11].g_word[7].r_bit.Q ;
  wire \g_bit[11].g_word[8].r_bit.Q ;
  wire \g_bit[11].g_word[9].r_bit.Q ;
  wire \g_bit[11].r_rs1.D ;
  wire \g_bit[11].r_rs1.Q ;
  wire \g_bit[11].r_rs2.D ;
  wire \g_bit[11].r_rs2.Q ;
  wire \g_bit[12].g_word[10].r_bit.Q ;
  wire \g_bit[12].g_word[11].r_bit.Q ;
  wire \g_bit[12].g_word[12].r_bit.Q ;
  wire \g_bit[12].g_word[13].r_bit.Q ;
  wire \g_bit[12].g_word[14].r_bit.Q ;
  wire \g_bit[12].g_word[15].r_bit.Q ;
  wire \g_bit[12].g_word[16].r_bit.Q ;
  wire \g_bit[12].g_word[17].r_bit.Q ;
  wire \g_bit[12].g_word[18].r_bit.Q ;
  wire \g_bit[12].g_word[19].r_bit.Q ;
  wire \g_bit[12].g_word[1].r_bit.Q ;
  wire \g_bit[12].g_word[20].r_bit.Q ;
  wire \g_bit[12].g_word[21].r_bit.Q ;
  wire \g_bit[12].g_word[22].r_bit.Q ;
  wire \g_bit[12].g_word[23].r_bit.Q ;
  wire \g_bit[12].g_word[24].r_bit.Q ;
  wire \g_bit[12].g_word[25].r_bit.Q ;
  wire \g_bit[12].g_word[26].r_bit.Q ;
  wire \g_bit[12].g_word[27].r_bit.Q ;
  wire \g_bit[12].g_word[28].r_bit.Q ;
  wire \g_bit[12].g_word[29].r_bit.Q ;
  wire \g_bit[12].g_word[2].r_bit.Q ;
  wire \g_bit[12].g_word[30].r_bit.Q ;
  wire \g_bit[12].g_word[31].r_bit.Q ;
  wire \g_bit[12].g_word[3].r_bit.Q ;
  wire \g_bit[12].g_word[4].r_bit.Q ;
  wire \g_bit[12].g_word[5].r_bit.Q ;
  wire \g_bit[12].g_word[6].r_bit.Q ;
  wire \g_bit[12].g_word[7].r_bit.Q ;
  wire \g_bit[12].g_word[8].r_bit.Q ;
  wire \g_bit[12].g_word[9].r_bit.Q ;
  wire \g_bit[12].r_rs1.D ;
  wire \g_bit[12].r_rs1.Q ;
  wire \g_bit[12].r_rs2.D ;
  wire \g_bit[12].r_rs2.Q ;
  wire \g_bit[13].g_word[10].r_bit.Q ;
  wire \g_bit[13].g_word[11].r_bit.Q ;
  wire \g_bit[13].g_word[12].r_bit.Q ;
  wire \g_bit[13].g_word[13].r_bit.Q ;
  wire \g_bit[13].g_word[14].r_bit.Q ;
  wire \g_bit[13].g_word[15].r_bit.Q ;
  wire \g_bit[13].g_word[16].r_bit.Q ;
  wire \g_bit[13].g_word[17].r_bit.Q ;
  wire \g_bit[13].g_word[18].r_bit.Q ;
  wire \g_bit[13].g_word[19].r_bit.Q ;
  wire \g_bit[13].g_word[1].r_bit.Q ;
  wire \g_bit[13].g_word[20].r_bit.Q ;
  wire \g_bit[13].g_word[21].r_bit.Q ;
  wire \g_bit[13].g_word[22].r_bit.Q ;
  wire \g_bit[13].g_word[23].r_bit.Q ;
  wire \g_bit[13].g_word[24].r_bit.Q ;
  wire \g_bit[13].g_word[25].r_bit.Q ;
  wire \g_bit[13].g_word[26].r_bit.Q ;
  wire \g_bit[13].g_word[27].r_bit.Q ;
  wire \g_bit[13].g_word[28].r_bit.Q ;
  wire \g_bit[13].g_word[29].r_bit.Q ;
  wire \g_bit[13].g_word[2].r_bit.Q ;
  wire \g_bit[13].g_word[30].r_bit.Q ;
  wire \g_bit[13].g_word[31].r_bit.Q ;
  wire \g_bit[13].g_word[3].r_bit.Q ;
  wire \g_bit[13].g_word[4].r_bit.Q ;
  wire \g_bit[13].g_word[5].r_bit.Q ;
  wire \g_bit[13].g_word[6].r_bit.Q ;
  wire \g_bit[13].g_word[7].r_bit.Q ;
  wire \g_bit[13].g_word[8].r_bit.Q ;
  wire \g_bit[13].g_word[9].r_bit.Q ;
  wire \g_bit[13].r_rs1.D ;
  wire \g_bit[13].r_rs1.Q ;
  wire \g_bit[13].r_rs2.D ;
  wire \g_bit[13].r_rs2.Q ;
  wire \g_bit[14].g_word[10].r_bit.Q ;
  wire \g_bit[14].g_word[11].r_bit.Q ;
  wire \g_bit[14].g_word[12].r_bit.Q ;
  wire \g_bit[14].g_word[13].r_bit.Q ;
  wire \g_bit[14].g_word[14].r_bit.Q ;
  wire \g_bit[14].g_word[15].r_bit.Q ;
  wire \g_bit[14].g_word[16].r_bit.Q ;
  wire \g_bit[14].g_word[17].r_bit.Q ;
  wire \g_bit[14].g_word[18].r_bit.Q ;
  wire \g_bit[14].g_word[19].r_bit.Q ;
  wire \g_bit[14].g_word[1].r_bit.Q ;
  wire \g_bit[14].g_word[20].r_bit.Q ;
  wire \g_bit[14].g_word[21].r_bit.Q ;
  wire \g_bit[14].g_word[22].r_bit.Q ;
  wire \g_bit[14].g_word[23].r_bit.Q ;
  wire \g_bit[14].g_word[24].r_bit.Q ;
  wire \g_bit[14].g_word[25].r_bit.Q ;
  wire \g_bit[14].g_word[26].r_bit.Q ;
  wire \g_bit[14].g_word[27].r_bit.Q ;
  wire \g_bit[14].g_word[28].r_bit.Q ;
  wire \g_bit[14].g_word[29].r_bit.Q ;
  wire \g_bit[14].g_word[2].r_bit.Q ;
  wire \g_bit[14].g_word[30].r_bit.Q ;
  wire \g_bit[14].g_word[31].r_bit.Q ;
  wire \g_bit[14].g_word[3].r_bit.Q ;
  wire \g_bit[14].g_word[4].r_bit.Q ;
  wire \g_bit[14].g_word[5].r_bit.Q ;
  wire \g_bit[14].g_word[6].r_bit.Q ;
  wire \g_bit[14].g_word[7].r_bit.Q ;
  wire \g_bit[14].g_word[8].r_bit.Q ;
  wire \g_bit[14].g_word[9].r_bit.Q ;
  wire \g_bit[14].r_rs1.D ;
  wire \g_bit[14].r_rs1.Q ;
  wire \g_bit[14].r_rs2.D ;
  wire \g_bit[14].r_rs2.Q ;
  wire \g_bit[15].g_word[10].r_bit.Q ;
  wire \g_bit[15].g_word[11].r_bit.Q ;
  wire \g_bit[15].g_word[12].r_bit.Q ;
  wire \g_bit[15].g_word[13].r_bit.Q ;
  wire \g_bit[15].g_word[14].r_bit.Q ;
  wire \g_bit[15].g_word[15].r_bit.Q ;
  wire \g_bit[15].g_word[16].r_bit.Q ;
  wire \g_bit[15].g_word[17].r_bit.Q ;
  wire \g_bit[15].g_word[18].r_bit.Q ;
  wire \g_bit[15].g_word[19].r_bit.Q ;
  wire \g_bit[15].g_word[1].r_bit.Q ;
  wire \g_bit[15].g_word[20].r_bit.Q ;
  wire \g_bit[15].g_word[21].r_bit.Q ;
  wire \g_bit[15].g_word[22].r_bit.Q ;
  wire \g_bit[15].g_word[23].r_bit.Q ;
  wire \g_bit[15].g_word[24].r_bit.Q ;
  wire \g_bit[15].g_word[25].r_bit.Q ;
  wire \g_bit[15].g_word[26].r_bit.Q ;
  wire \g_bit[15].g_word[27].r_bit.Q ;
  wire \g_bit[15].g_word[28].r_bit.Q ;
  wire \g_bit[15].g_word[29].r_bit.Q ;
  wire \g_bit[15].g_word[2].r_bit.Q ;
  wire \g_bit[15].g_word[30].r_bit.Q ;
  wire \g_bit[15].g_word[31].r_bit.Q ;
  wire \g_bit[15].g_word[3].r_bit.Q ;
  wire \g_bit[15].g_word[4].r_bit.Q ;
  wire \g_bit[15].g_word[5].r_bit.Q ;
  wire \g_bit[15].g_word[6].r_bit.Q ;
  wire \g_bit[15].g_word[7].r_bit.Q ;
  wire \g_bit[15].g_word[8].r_bit.Q ;
  wire \g_bit[15].g_word[9].r_bit.Q ;
  wire \g_bit[15].r_rs1.D ;
  wire \g_bit[15].r_rs1.Q ;
  wire \g_bit[15].r_rs2.D ;
  wire \g_bit[15].r_rs2.Q ;
  wire \g_bit[16].g_word[10].r_bit.Q ;
  wire \g_bit[16].g_word[11].r_bit.Q ;
  wire \g_bit[16].g_word[12].r_bit.Q ;
  wire \g_bit[16].g_word[13].r_bit.Q ;
  wire \g_bit[16].g_word[14].r_bit.Q ;
  wire \g_bit[16].g_word[15].r_bit.Q ;
  wire \g_bit[16].g_word[16].r_bit.Q ;
  wire \g_bit[16].g_word[17].r_bit.Q ;
  wire \g_bit[16].g_word[18].r_bit.Q ;
  wire \g_bit[16].g_word[19].r_bit.Q ;
  wire \g_bit[16].g_word[1].r_bit.Q ;
  wire \g_bit[16].g_word[20].r_bit.Q ;
  wire \g_bit[16].g_word[21].r_bit.Q ;
  wire \g_bit[16].g_word[22].r_bit.Q ;
  wire \g_bit[16].g_word[23].r_bit.Q ;
  wire \g_bit[16].g_word[24].r_bit.Q ;
  wire \g_bit[16].g_word[25].r_bit.Q ;
  wire \g_bit[16].g_word[26].r_bit.Q ;
  wire \g_bit[16].g_word[27].r_bit.Q ;
  wire \g_bit[16].g_word[28].r_bit.Q ;
  wire \g_bit[16].g_word[29].r_bit.Q ;
  wire \g_bit[16].g_word[2].r_bit.Q ;
  wire \g_bit[16].g_word[30].r_bit.Q ;
  wire \g_bit[16].g_word[31].r_bit.Q ;
  wire \g_bit[16].g_word[3].r_bit.Q ;
  wire \g_bit[16].g_word[4].r_bit.Q ;
  wire \g_bit[16].g_word[5].r_bit.Q ;
  wire \g_bit[16].g_word[6].r_bit.Q ;
  wire \g_bit[16].g_word[7].r_bit.Q ;
  wire \g_bit[16].g_word[8].r_bit.Q ;
  wire \g_bit[16].g_word[9].r_bit.Q ;
  wire \g_bit[16].r_rs1.D ;
  wire \g_bit[16].r_rs1.Q ;
  wire \g_bit[16].r_rs2.D ;
  wire \g_bit[16].r_rs2.Q ;
  wire \g_bit[17].g_word[10].r_bit.Q ;
  wire \g_bit[17].g_word[11].r_bit.Q ;
  wire \g_bit[17].g_word[12].r_bit.Q ;
  wire \g_bit[17].g_word[13].r_bit.Q ;
  wire \g_bit[17].g_word[14].r_bit.Q ;
  wire \g_bit[17].g_word[15].r_bit.Q ;
  wire \g_bit[17].g_word[16].r_bit.Q ;
  wire \g_bit[17].g_word[17].r_bit.Q ;
  wire \g_bit[17].g_word[18].r_bit.Q ;
  wire \g_bit[17].g_word[19].r_bit.Q ;
  wire \g_bit[17].g_word[1].r_bit.Q ;
  wire \g_bit[17].g_word[20].r_bit.Q ;
  wire \g_bit[17].g_word[21].r_bit.Q ;
  wire \g_bit[17].g_word[22].r_bit.Q ;
  wire \g_bit[17].g_word[23].r_bit.Q ;
  wire \g_bit[17].g_word[24].r_bit.Q ;
  wire \g_bit[17].g_word[25].r_bit.Q ;
  wire \g_bit[17].g_word[26].r_bit.Q ;
  wire \g_bit[17].g_word[27].r_bit.Q ;
  wire \g_bit[17].g_word[28].r_bit.Q ;
  wire \g_bit[17].g_word[29].r_bit.Q ;
  wire \g_bit[17].g_word[2].r_bit.Q ;
  wire \g_bit[17].g_word[30].r_bit.Q ;
  wire \g_bit[17].g_word[31].r_bit.Q ;
  wire \g_bit[17].g_word[3].r_bit.Q ;
  wire \g_bit[17].g_word[4].r_bit.Q ;
  wire \g_bit[17].g_word[5].r_bit.Q ;
  wire \g_bit[17].g_word[6].r_bit.Q ;
  wire \g_bit[17].g_word[7].r_bit.Q ;
  wire \g_bit[17].g_word[8].r_bit.Q ;
  wire \g_bit[17].g_word[9].r_bit.Q ;
  wire \g_bit[17].r_rs1.D ;
  wire \g_bit[17].r_rs1.Q ;
  wire \g_bit[17].r_rs2.D ;
  wire \g_bit[17].r_rs2.Q ;
  wire \g_bit[18].g_word[10].r_bit.Q ;
  wire \g_bit[18].g_word[11].r_bit.Q ;
  wire \g_bit[18].g_word[12].r_bit.Q ;
  wire \g_bit[18].g_word[13].r_bit.Q ;
  wire \g_bit[18].g_word[14].r_bit.Q ;
  wire \g_bit[18].g_word[15].r_bit.Q ;
  wire \g_bit[18].g_word[16].r_bit.Q ;
  wire \g_bit[18].g_word[17].r_bit.Q ;
  wire \g_bit[18].g_word[18].r_bit.Q ;
  wire \g_bit[18].g_word[19].r_bit.Q ;
  wire \g_bit[18].g_word[1].r_bit.Q ;
  wire \g_bit[18].g_word[20].r_bit.Q ;
  wire \g_bit[18].g_word[21].r_bit.Q ;
  wire \g_bit[18].g_word[22].r_bit.Q ;
  wire \g_bit[18].g_word[23].r_bit.Q ;
  wire \g_bit[18].g_word[24].r_bit.Q ;
  wire \g_bit[18].g_word[25].r_bit.Q ;
  wire \g_bit[18].g_word[26].r_bit.Q ;
  wire \g_bit[18].g_word[27].r_bit.Q ;
  wire \g_bit[18].g_word[28].r_bit.Q ;
  wire \g_bit[18].g_word[29].r_bit.Q ;
  wire \g_bit[18].g_word[2].r_bit.Q ;
  wire \g_bit[18].g_word[30].r_bit.Q ;
  wire \g_bit[18].g_word[31].r_bit.Q ;
  wire \g_bit[18].g_word[3].r_bit.Q ;
  wire \g_bit[18].g_word[4].r_bit.Q ;
  wire \g_bit[18].g_word[5].r_bit.Q ;
  wire \g_bit[18].g_word[6].r_bit.Q ;
  wire \g_bit[18].g_word[7].r_bit.Q ;
  wire \g_bit[18].g_word[8].r_bit.Q ;
  wire \g_bit[18].g_word[9].r_bit.Q ;
  wire \g_bit[18].r_rs1.D ;
  wire \g_bit[18].r_rs1.Q ;
  wire \g_bit[18].r_rs2.D ;
  wire \g_bit[18].r_rs2.Q ;
  wire \g_bit[19].g_word[10].r_bit.Q ;
  wire \g_bit[19].g_word[11].r_bit.Q ;
  wire \g_bit[19].g_word[12].r_bit.Q ;
  wire \g_bit[19].g_word[13].r_bit.Q ;
  wire \g_bit[19].g_word[14].r_bit.Q ;
  wire \g_bit[19].g_word[15].r_bit.Q ;
  wire \g_bit[19].g_word[16].r_bit.Q ;
  wire \g_bit[19].g_word[17].r_bit.Q ;
  wire \g_bit[19].g_word[18].r_bit.Q ;
  wire \g_bit[19].g_word[19].r_bit.Q ;
  wire \g_bit[19].g_word[1].r_bit.Q ;
  wire \g_bit[19].g_word[20].r_bit.Q ;
  wire \g_bit[19].g_word[21].r_bit.Q ;
  wire \g_bit[19].g_word[22].r_bit.Q ;
  wire \g_bit[19].g_word[23].r_bit.Q ;
  wire \g_bit[19].g_word[24].r_bit.Q ;
  wire \g_bit[19].g_word[25].r_bit.Q ;
  wire \g_bit[19].g_word[26].r_bit.Q ;
  wire \g_bit[19].g_word[27].r_bit.Q ;
  wire \g_bit[19].g_word[28].r_bit.Q ;
  wire \g_bit[19].g_word[29].r_bit.Q ;
  wire \g_bit[19].g_word[2].r_bit.Q ;
  wire \g_bit[19].g_word[30].r_bit.Q ;
  wire \g_bit[19].g_word[31].r_bit.Q ;
  wire \g_bit[19].g_word[3].r_bit.Q ;
  wire \g_bit[19].g_word[4].r_bit.Q ;
  wire \g_bit[19].g_word[5].r_bit.Q ;
  wire \g_bit[19].g_word[6].r_bit.Q ;
  wire \g_bit[19].g_word[7].r_bit.Q ;
  wire \g_bit[19].g_word[8].r_bit.Q ;
  wire \g_bit[19].g_word[9].r_bit.Q ;
  wire \g_bit[19].r_rs1.D ;
  wire \g_bit[19].r_rs1.Q ;
  wire \g_bit[19].r_rs2.D ;
  wire \g_bit[19].r_rs2.Q ;
  wire \g_bit[1].g_word[10].r_bit.Q ;
  wire \g_bit[1].g_word[11].r_bit.Q ;
  wire \g_bit[1].g_word[12].r_bit.Q ;
  wire \g_bit[1].g_word[13].r_bit.Q ;
  wire \g_bit[1].g_word[14].r_bit.Q ;
  wire \g_bit[1].g_word[15].r_bit.Q ;
  wire \g_bit[1].g_word[16].r_bit.Q ;
  wire \g_bit[1].g_word[17].r_bit.Q ;
  wire \g_bit[1].g_word[18].r_bit.Q ;
  wire \g_bit[1].g_word[19].r_bit.Q ;
  wire \g_bit[1].g_word[1].r_bit.Q ;
  wire \g_bit[1].g_word[20].r_bit.Q ;
  wire \g_bit[1].g_word[21].r_bit.Q ;
  wire \g_bit[1].g_word[22].r_bit.Q ;
  wire \g_bit[1].g_word[23].r_bit.Q ;
  wire \g_bit[1].g_word[24].r_bit.Q ;
  wire \g_bit[1].g_word[25].r_bit.Q ;
  wire \g_bit[1].g_word[26].r_bit.Q ;
  wire \g_bit[1].g_word[27].r_bit.Q ;
  wire \g_bit[1].g_word[28].r_bit.Q ;
  wire \g_bit[1].g_word[29].r_bit.Q ;
  wire \g_bit[1].g_word[2].r_bit.Q ;
  wire \g_bit[1].g_word[30].r_bit.Q ;
  wire \g_bit[1].g_word[31].r_bit.Q ;
  wire \g_bit[1].g_word[3].r_bit.Q ;
  wire \g_bit[1].g_word[4].r_bit.Q ;
  wire \g_bit[1].g_word[5].r_bit.Q ;
  wire \g_bit[1].g_word[6].r_bit.Q ;
  wire \g_bit[1].g_word[7].r_bit.Q ;
  wire \g_bit[1].g_word[8].r_bit.Q ;
  wire \g_bit[1].g_word[9].r_bit.Q ;
  wire \g_bit[1].r_rs1.D ;
  wire \g_bit[1].r_rs1.Q ;
  wire \g_bit[1].r_rs2.D ;
  wire \g_bit[1].r_rs2.Q ;
  wire \g_bit[20].g_word[10].r_bit.Q ;
  wire \g_bit[20].g_word[11].r_bit.Q ;
  wire \g_bit[20].g_word[12].r_bit.Q ;
  wire \g_bit[20].g_word[13].r_bit.Q ;
  wire \g_bit[20].g_word[14].r_bit.Q ;
  wire \g_bit[20].g_word[15].r_bit.Q ;
  wire \g_bit[20].g_word[16].r_bit.Q ;
  wire \g_bit[20].g_word[17].r_bit.Q ;
  wire \g_bit[20].g_word[18].r_bit.Q ;
  wire \g_bit[20].g_word[19].r_bit.Q ;
  wire \g_bit[20].g_word[1].r_bit.Q ;
  wire \g_bit[20].g_word[20].r_bit.Q ;
  wire \g_bit[20].g_word[21].r_bit.Q ;
  wire \g_bit[20].g_word[22].r_bit.Q ;
  wire \g_bit[20].g_word[23].r_bit.Q ;
  wire \g_bit[20].g_word[24].r_bit.Q ;
  wire \g_bit[20].g_word[25].r_bit.Q ;
  wire \g_bit[20].g_word[26].r_bit.Q ;
  wire \g_bit[20].g_word[27].r_bit.Q ;
  wire \g_bit[20].g_word[28].r_bit.Q ;
  wire \g_bit[20].g_word[29].r_bit.Q ;
  wire \g_bit[20].g_word[2].r_bit.Q ;
  wire \g_bit[20].g_word[30].r_bit.Q ;
  wire \g_bit[20].g_word[31].r_bit.Q ;
  wire \g_bit[20].g_word[3].r_bit.Q ;
  wire \g_bit[20].g_word[4].r_bit.Q ;
  wire \g_bit[20].g_word[5].r_bit.Q ;
  wire \g_bit[20].g_word[6].r_bit.Q ;
  wire \g_bit[20].g_word[7].r_bit.Q ;
  wire \g_bit[20].g_word[8].r_bit.Q ;
  wire \g_bit[20].g_word[9].r_bit.Q ;
  wire \g_bit[20].r_rs1.D ;
  wire \g_bit[20].r_rs1.Q ;
  wire \g_bit[20].r_rs2.D ;
  wire \g_bit[20].r_rs2.Q ;
  wire \g_bit[21].g_word[10].r_bit.Q ;
  wire \g_bit[21].g_word[11].r_bit.Q ;
  wire \g_bit[21].g_word[12].r_bit.Q ;
  wire \g_bit[21].g_word[13].r_bit.Q ;
  wire \g_bit[21].g_word[14].r_bit.Q ;
  wire \g_bit[21].g_word[15].r_bit.Q ;
  wire \g_bit[21].g_word[16].r_bit.Q ;
  wire \g_bit[21].g_word[17].r_bit.Q ;
  wire \g_bit[21].g_word[18].r_bit.Q ;
  wire \g_bit[21].g_word[19].r_bit.Q ;
  wire \g_bit[21].g_word[1].r_bit.Q ;
  wire \g_bit[21].g_word[20].r_bit.Q ;
  wire \g_bit[21].g_word[21].r_bit.Q ;
  wire \g_bit[21].g_word[22].r_bit.Q ;
  wire \g_bit[21].g_word[23].r_bit.Q ;
  wire \g_bit[21].g_word[24].r_bit.Q ;
  wire \g_bit[21].g_word[25].r_bit.Q ;
  wire \g_bit[21].g_word[26].r_bit.Q ;
  wire \g_bit[21].g_word[27].r_bit.Q ;
  wire \g_bit[21].g_word[28].r_bit.Q ;
  wire \g_bit[21].g_word[29].r_bit.Q ;
  wire \g_bit[21].g_word[2].r_bit.Q ;
  wire \g_bit[21].g_word[30].r_bit.Q ;
  wire \g_bit[21].g_word[31].r_bit.Q ;
  wire \g_bit[21].g_word[3].r_bit.Q ;
  wire \g_bit[21].g_word[4].r_bit.Q ;
  wire \g_bit[21].g_word[5].r_bit.Q ;
  wire \g_bit[21].g_word[6].r_bit.Q ;
  wire \g_bit[21].g_word[7].r_bit.Q ;
  wire \g_bit[21].g_word[8].r_bit.Q ;
  wire \g_bit[21].g_word[9].r_bit.Q ;
  wire \g_bit[21].r_rs1.D ;
  wire \g_bit[21].r_rs1.Q ;
  wire \g_bit[21].r_rs2.D ;
  wire \g_bit[21].r_rs2.Q ;
  wire \g_bit[22].g_word[10].r_bit.Q ;
  wire \g_bit[22].g_word[11].r_bit.Q ;
  wire \g_bit[22].g_word[12].r_bit.Q ;
  wire \g_bit[22].g_word[13].r_bit.Q ;
  wire \g_bit[22].g_word[14].r_bit.Q ;
  wire \g_bit[22].g_word[15].r_bit.Q ;
  wire \g_bit[22].g_word[16].r_bit.Q ;
  wire \g_bit[22].g_word[17].r_bit.Q ;
  wire \g_bit[22].g_word[18].r_bit.Q ;
  wire \g_bit[22].g_word[19].r_bit.Q ;
  wire \g_bit[22].g_word[1].r_bit.Q ;
  wire \g_bit[22].g_word[20].r_bit.Q ;
  wire \g_bit[22].g_word[21].r_bit.Q ;
  wire \g_bit[22].g_word[22].r_bit.Q ;
  wire \g_bit[22].g_word[23].r_bit.Q ;
  wire \g_bit[22].g_word[24].r_bit.Q ;
  wire \g_bit[22].g_word[25].r_bit.Q ;
  wire \g_bit[22].g_word[26].r_bit.Q ;
  wire \g_bit[22].g_word[27].r_bit.Q ;
  wire \g_bit[22].g_word[28].r_bit.Q ;
  wire \g_bit[22].g_word[29].r_bit.Q ;
  wire \g_bit[22].g_word[2].r_bit.Q ;
  wire \g_bit[22].g_word[30].r_bit.Q ;
  wire \g_bit[22].g_word[31].r_bit.Q ;
  wire \g_bit[22].g_word[3].r_bit.Q ;
  wire \g_bit[22].g_word[4].r_bit.Q ;
  wire \g_bit[22].g_word[5].r_bit.Q ;
  wire \g_bit[22].g_word[6].r_bit.Q ;
  wire \g_bit[22].g_word[7].r_bit.Q ;
  wire \g_bit[22].g_word[8].r_bit.Q ;
  wire \g_bit[22].g_word[9].r_bit.Q ;
  wire \g_bit[22].r_rs1.D ;
  wire \g_bit[22].r_rs1.Q ;
  wire \g_bit[22].r_rs2.D ;
  wire \g_bit[22].r_rs2.Q ;
  wire \g_bit[23].g_word[10].r_bit.Q ;
  wire \g_bit[23].g_word[11].r_bit.Q ;
  wire \g_bit[23].g_word[12].r_bit.Q ;
  wire \g_bit[23].g_word[13].r_bit.Q ;
  wire \g_bit[23].g_word[14].r_bit.Q ;
  wire \g_bit[23].g_word[15].r_bit.Q ;
  wire \g_bit[23].g_word[16].r_bit.Q ;
  wire \g_bit[23].g_word[17].r_bit.Q ;
  wire \g_bit[23].g_word[18].r_bit.Q ;
  wire \g_bit[23].g_word[19].r_bit.Q ;
  wire \g_bit[23].g_word[1].r_bit.Q ;
  wire \g_bit[23].g_word[20].r_bit.Q ;
  wire \g_bit[23].g_word[21].r_bit.Q ;
  wire \g_bit[23].g_word[22].r_bit.Q ;
  wire \g_bit[23].g_word[23].r_bit.Q ;
  wire \g_bit[23].g_word[24].r_bit.Q ;
  wire \g_bit[23].g_word[25].r_bit.Q ;
  wire \g_bit[23].g_word[26].r_bit.Q ;
  wire \g_bit[23].g_word[27].r_bit.Q ;
  wire \g_bit[23].g_word[28].r_bit.Q ;
  wire \g_bit[23].g_word[29].r_bit.Q ;
  wire \g_bit[23].g_word[2].r_bit.Q ;
  wire \g_bit[23].g_word[30].r_bit.Q ;
  wire \g_bit[23].g_word[31].r_bit.Q ;
  wire \g_bit[23].g_word[3].r_bit.Q ;
  wire \g_bit[23].g_word[4].r_bit.Q ;
  wire \g_bit[23].g_word[5].r_bit.Q ;
  wire \g_bit[23].g_word[6].r_bit.Q ;
  wire \g_bit[23].g_word[7].r_bit.Q ;
  wire \g_bit[23].g_word[8].r_bit.Q ;
  wire \g_bit[23].g_word[9].r_bit.Q ;
  wire \g_bit[23].r_rs1.D ;
  wire \g_bit[23].r_rs1.Q ;
  wire \g_bit[23].r_rs2.D ;
  wire \g_bit[23].r_rs2.Q ;
  wire \g_bit[24].g_word[10].r_bit.Q ;
  wire \g_bit[24].g_word[11].r_bit.Q ;
  wire \g_bit[24].g_word[12].r_bit.Q ;
  wire \g_bit[24].g_word[13].r_bit.Q ;
  wire \g_bit[24].g_word[14].r_bit.Q ;
  wire \g_bit[24].g_word[15].r_bit.Q ;
  wire \g_bit[24].g_word[16].r_bit.Q ;
  wire \g_bit[24].g_word[17].r_bit.Q ;
  wire \g_bit[24].g_word[18].r_bit.Q ;
  wire \g_bit[24].g_word[19].r_bit.Q ;
  wire \g_bit[24].g_word[1].r_bit.Q ;
  wire \g_bit[24].g_word[20].r_bit.Q ;
  wire \g_bit[24].g_word[21].r_bit.Q ;
  wire \g_bit[24].g_word[22].r_bit.Q ;
  wire \g_bit[24].g_word[23].r_bit.Q ;
  wire \g_bit[24].g_word[24].r_bit.Q ;
  wire \g_bit[24].g_word[25].r_bit.Q ;
  wire \g_bit[24].g_word[26].r_bit.Q ;
  wire \g_bit[24].g_word[27].r_bit.Q ;
  wire \g_bit[24].g_word[28].r_bit.Q ;
  wire \g_bit[24].g_word[29].r_bit.Q ;
  wire \g_bit[24].g_word[2].r_bit.Q ;
  wire \g_bit[24].g_word[30].r_bit.Q ;
  wire \g_bit[24].g_word[31].r_bit.Q ;
  wire \g_bit[24].g_word[3].r_bit.Q ;
  wire \g_bit[24].g_word[4].r_bit.Q ;
  wire \g_bit[24].g_word[5].r_bit.Q ;
  wire \g_bit[24].g_word[6].r_bit.Q ;
  wire \g_bit[24].g_word[7].r_bit.Q ;
  wire \g_bit[24].g_word[8].r_bit.Q ;
  wire \g_bit[24].g_word[9].r_bit.Q ;
  wire \g_bit[24].r_rs1.D ;
  wire \g_bit[24].r_rs1.Q ;
  wire \g_bit[24].r_rs2.D ;
  wire \g_bit[24].r_rs2.Q ;
  wire \g_bit[25].g_word[10].r_bit.Q ;
  wire \g_bit[25].g_word[11].r_bit.Q ;
  wire \g_bit[25].g_word[12].r_bit.Q ;
  wire \g_bit[25].g_word[13].r_bit.Q ;
  wire \g_bit[25].g_word[14].r_bit.Q ;
  wire \g_bit[25].g_word[15].r_bit.Q ;
  wire \g_bit[25].g_word[16].r_bit.Q ;
  wire \g_bit[25].g_word[17].r_bit.Q ;
  wire \g_bit[25].g_word[18].r_bit.Q ;
  wire \g_bit[25].g_word[19].r_bit.Q ;
  wire \g_bit[25].g_word[1].r_bit.Q ;
  wire \g_bit[25].g_word[20].r_bit.Q ;
  wire \g_bit[25].g_word[21].r_bit.Q ;
  wire \g_bit[25].g_word[22].r_bit.Q ;
  wire \g_bit[25].g_word[23].r_bit.Q ;
  wire \g_bit[25].g_word[24].r_bit.Q ;
  wire \g_bit[25].g_word[25].r_bit.Q ;
  wire \g_bit[25].g_word[26].r_bit.Q ;
  wire \g_bit[25].g_word[27].r_bit.Q ;
  wire \g_bit[25].g_word[28].r_bit.Q ;
  wire \g_bit[25].g_word[29].r_bit.Q ;
  wire \g_bit[25].g_word[2].r_bit.Q ;
  wire \g_bit[25].g_word[30].r_bit.Q ;
  wire \g_bit[25].g_word[31].r_bit.Q ;
  wire \g_bit[25].g_word[3].r_bit.Q ;
  wire \g_bit[25].g_word[4].r_bit.Q ;
  wire \g_bit[25].g_word[5].r_bit.Q ;
  wire \g_bit[25].g_word[6].r_bit.Q ;
  wire \g_bit[25].g_word[7].r_bit.Q ;
  wire \g_bit[25].g_word[8].r_bit.Q ;
  wire \g_bit[25].g_word[9].r_bit.Q ;
  wire \g_bit[25].r_rs1.D ;
  wire \g_bit[25].r_rs1.Q ;
  wire \g_bit[25].r_rs2.D ;
  wire \g_bit[25].r_rs2.Q ;
  wire \g_bit[26].g_word[10].r_bit.Q ;
  wire \g_bit[26].g_word[11].r_bit.Q ;
  wire \g_bit[26].g_word[12].r_bit.Q ;
  wire \g_bit[26].g_word[13].r_bit.Q ;
  wire \g_bit[26].g_word[14].r_bit.Q ;
  wire \g_bit[26].g_word[15].r_bit.Q ;
  wire \g_bit[26].g_word[16].r_bit.Q ;
  wire \g_bit[26].g_word[17].r_bit.Q ;
  wire \g_bit[26].g_word[18].r_bit.Q ;
  wire \g_bit[26].g_word[19].r_bit.Q ;
  wire \g_bit[26].g_word[1].r_bit.Q ;
  wire \g_bit[26].g_word[20].r_bit.Q ;
  wire \g_bit[26].g_word[21].r_bit.Q ;
  wire \g_bit[26].g_word[22].r_bit.Q ;
  wire \g_bit[26].g_word[23].r_bit.Q ;
  wire \g_bit[26].g_word[24].r_bit.Q ;
  wire \g_bit[26].g_word[25].r_bit.Q ;
  wire \g_bit[26].g_word[26].r_bit.Q ;
  wire \g_bit[26].g_word[27].r_bit.Q ;
  wire \g_bit[26].g_word[28].r_bit.Q ;
  wire \g_bit[26].g_word[29].r_bit.Q ;
  wire \g_bit[26].g_word[2].r_bit.Q ;
  wire \g_bit[26].g_word[30].r_bit.Q ;
  wire \g_bit[26].g_word[31].r_bit.Q ;
  wire \g_bit[26].g_word[3].r_bit.Q ;
  wire \g_bit[26].g_word[4].r_bit.Q ;
  wire \g_bit[26].g_word[5].r_bit.Q ;
  wire \g_bit[26].g_word[6].r_bit.Q ;
  wire \g_bit[26].g_word[7].r_bit.Q ;
  wire \g_bit[26].g_word[8].r_bit.Q ;
  wire \g_bit[26].g_word[9].r_bit.Q ;
  wire \g_bit[26].r_rs1.D ;
  wire \g_bit[26].r_rs1.Q ;
  wire \g_bit[26].r_rs2.D ;
  wire \g_bit[26].r_rs2.Q ;
  wire \g_bit[27].g_word[10].r_bit.Q ;
  wire \g_bit[27].g_word[11].r_bit.Q ;
  wire \g_bit[27].g_word[12].r_bit.Q ;
  wire \g_bit[27].g_word[13].r_bit.Q ;
  wire \g_bit[27].g_word[14].r_bit.Q ;
  wire \g_bit[27].g_word[15].r_bit.Q ;
  wire \g_bit[27].g_word[16].r_bit.Q ;
  wire \g_bit[27].g_word[17].r_bit.Q ;
  wire \g_bit[27].g_word[18].r_bit.Q ;
  wire \g_bit[27].g_word[19].r_bit.Q ;
  wire \g_bit[27].g_word[1].r_bit.Q ;
  wire \g_bit[27].g_word[20].r_bit.Q ;
  wire \g_bit[27].g_word[21].r_bit.Q ;
  wire \g_bit[27].g_word[22].r_bit.Q ;
  wire \g_bit[27].g_word[23].r_bit.Q ;
  wire \g_bit[27].g_word[24].r_bit.Q ;
  wire \g_bit[27].g_word[25].r_bit.Q ;
  wire \g_bit[27].g_word[26].r_bit.Q ;
  wire \g_bit[27].g_word[27].r_bit.Q ;
  wire \g_bit[27].g_word[28].r_bit.Q ;
  wire \g_bit[27].g_word[29].r_bit.Q ;
  wire \g_bit[27].g_word[2].r_bit.Q ;
  wire \g_bit[27].g_word[30].r_bit.Q ;
  wire \g_bit[27].g_word[31].r_bit.Q ;
  wire \g_bit[27].g_word[3].r_bit.Q ;
  wire \g_bit[27].g_word[4].r_bit.Q ;
  wire \g_bit[27].g_word[5].r_bit.Q ;
  wire \g_bit[27].g_word[6].r_bit.Q ;
  wire \g_bit[27].g_word[7].r_bit.Q ;
  wire \g_bit[27].g_word[8].r_bit.Q ;
  wire \g_bit[27].g_word[9].r_bit.Q ;
  wire \g_bit[27].r_rs1.D ;
  wire \g_bit[27].r_rs1.Q ;
  wire \g_bit[27].r_rs2.D ;
  wire \g_bit[27].r_rs2.Q ;
  wire \g_bit[28].g_word[10].r_bit.Q ;
  wire \g_bit[28].g_word[11].r_bit.Q ;
  wire \g_bit[28].g_word[12].r_bit.Q ;
  wire \g_bit[28].g_word[13].r_bit.Q ;
  wire \g_bit[28].g_word[14].r_bit.Q ;
  wire \g_bit[28].g_word[15].r_bit.Q ;
  wire \g_bit[28].g_word[16].r_bit.Q ;
  wire \g_bit[28].g_word[17].r_bit.Q ;
  wire \g_bit[28].g_word[18].r_bit.Q ;
  wire \g_bit[28].g_word[19].r_bit.Q ;
  wire \g_bit[28].g_word[1].r_bit.Q ;
  wire \g_bit[28].g_word[20].r_bit.Q ;
  wire \g_bit[28].g_word[21].r_bit.Q ;
  wire \g_bit[28].g_word[22].r_bit.Q ;
  wire \g_bit[28].g_word[23].r_bit.Q ;
  wire \g_bit[28].g_word[24].r_bit.Q ;
  wire \g_bit[28].g_word[25].r_bit.Q ;
  wire \g_bit[28].g_word[26].r_bit.Q ;
  wire \g_bit[28].g_word[27].r_bit.Q ;
  wire \g_bit[28].g_word[28].r_bit.Q ;
  wire \g_bit[28].g_word[29].r_bit.Q ;
  wire \g_bit[28].g_word[2].r_bit.Q ;
  wire \g_bit[28].g_word[30].r_bit.Q ;
  wire \g_bit[28].g_word[31].r_bit.Q ;
  wire \g_bit[28].g_word[3].r_bit.Q ;
  wire \g_bit[28].g_word[4].r_bit.Q ;
  wire \g_bit[28].g_word[5].r_bit.Q ;
  wire \g_bit[28].g_word[6].r_bit.Q ;
  wire \g_bit[28].g_word[7].r_bit.Q ;
  wire \g_bit[28].g_word[8].r_bit.Q ;
  wire \g_bit[28].g_word[9].r_bit.Q ;
  wire \g_bit[28].r_rs1.D ;
  wire \g_bit[28].r_rs1.Q ;
  wire \g_bit[28].r_rs2.D ;
  wire \g_bit[28].r_rs2.Q ;
  wire \g_bit[29].g_word[10].r_bit.Q ;
  wire \g_bit[29].g_word[11].r_bit.Q ;
  wire \g_bit[29].g_word[12].r_bit.Q ;
  wire \g_bit[29].g_word[13].r_bit.Q ;
  wire \g_bit[29].g_word[14].r_bit.Q ;
  wire \g_bit[29].g_word[15].r_bit.Q ;
  wire \g_bit[29].g_word[16].r_bit.Q ;
  wire \g_bit[29].g_word[17].r_bit.Q ;
  wire \g_bit[29].g_word[18].r_bit.Q ;
  wire \g_bit[29].g_word[19].r_bit.Q ;
  wire \g_bit[29].g_word[1].r_bit.Q ;
  wire \g_bit[29].g_word[20].r_bit.Q ;
  wire \g_bit[29].g_word[21].r_bit.Q ;
  wire \g_bit[29].g_word[22].r_bit.Q ;
  wire \g_bit[29].g_word[23].r_bit.Q ;
  wire \g_bit[29].g_word[24].r_bit.Q ;
  wire \g_bit[29].g_word[25].r_bit.Q ;
  wire \g_bit[29].g_word[26].r_bit.Q ;
  wire \g_bit[29].g_word[27].r_bit.Q ;
  wire \g_bit[29].g_word[28].r_bit.Q ;
  wire \g_bit[29].g_word[29].r_bit.Q ;
  wire \g_bit[29].g_word[2].r_bit.Q ;
  wire \g_bit[29].g_word[30].r_bit.Q ;
  wire \g_bit[29].g_word[31].r_bit.Q ;
  wire \g_bit[29].g_word[3].r_bit.Q ;
  wire \g_bit[29].g_word[4].r_bit.Q ;
  wire \g_bit[29].g_word[5].r_bit.Q ;
  wire \g_bit[29].g_word[6].r_bit.Q ;
  wire \g_bit[29].g_word[7].r_bit.Q ;
  wire \g_bit[29].g_word[8].r_bit.Q ;
  wire \g_bit[29].g_word[9].r_bit.Q ;
  wire \g_bit[29].r_rs1.D ;
  wire \g_bit[29].r_rs1.Q ;
  wire \g_bit[29].r_rs2.D ;
  wire \g_bit[29].r_rs2.Q ;
  wire \g_bit[2].g_word[10].r_bit.Q ;
  wire \g_bit[2].g_word[11].r_bit.Q ;
  wire \g_bit[2].g_word[12].r_bit.Q ;
  wire \g_bit[2].g_word[13].r_bit.Q ;
  wire \g_bit[2].g_word[14].r_bit.Q ;
  wire \g_bit[2].g_word[15].r_bit.Q ;
  wire \g_bit[2].g_word[16].r_bit.Q ;
  wire \g_bit[2].g_word[17].r_bit.Q ;
  wire \g_bit[2].g_word[18].r_bit.Q ;
  wire \g_bit[2].g_word[19].r_bit.Q ;
  wire \g_bit[2].g_word[1].r_bit.Q ;
  wire \g_bit[2].g_word[20].r_bit.Q ;
  wire \g_bit[2].g_word[21].r_bit.Q ;
  wire \g_bit[2].g_word[22].r_bit.Q ;
  wire \g_bit[2].g_word[23].r_bit.Q ;
  wire \g_bit[2].g_word[24].r_bit.Q ;
  wire \g_bit[2].g_word[25].r_bit.Q ;
  wire \g_bit[2].g_word[26].r_bit.Q ;
  wire \g_bit[2].g_word[27].r_bit.Q ;
  wire \g_bit[2].g_word[28].r_bit.Q ;
  wire \g_bit[2].g_word[29].r_bit.Q ;
  wire \g_bit[2].g_word[2].r_bit.Q ;
  wire \g_bit[2].g_word[30].r_bit.Q ;
  wire \g_bit[2].g_word[31].r_bit.Q ;
  wire \g_bit[2].g_word[3].r_bit.Q ;
  wire \g_bit[2].g_word[4].r_bit.Q ;
  wire \g_bit[2].g_word[5].r_bit.Q ;
  wire \g_bit[2].g_word[6].r_bit.Q ;
  wire \g_bit[2].g_word[7].r_bit.Q ;
  wire \g_bit[2].g_word[8].r_bit.Q ;
  wire \g_bit[2].g_word[9].r_bit.Q ;
  wire \g_bit[2].r_rs1.D ;
  wire \g_bit[2].r_rs1.Q ;
  wire \g_bit[2].r_rs2.D ;
  wire \g_bit[2].r_rs2.Q ;
  wire \g_bit[30].g_word[10].r_bit.Q ;
  wire \g_bit[30].g_word[11].r_bit.Q ;
  wire \g_bit[30].g_word[12].r_bit.Q ;
  wire \g_bit[30].g_word[13].r_bit.Q ;
  wire \g_bit[30].g_word[14].r_bit.Q ;
  wire \g_bit[30].g_word[15].r_bit.Q ;
  wire \g_bit[30].g_word[16].r_bit.Q ;
  wire \g_bit[30].g_word[17].r_bit.Q ;
  wire \g_bit[30].g_word[18].r_bit.Q ;
  wire \g_bit[30].g_word[19].r_bit.Q ;
  wire \g_bit[30].g_word[1].r_bit.Q ;
  wire \g_bit[30].g_word[20].r_bit.Q ;
  wire \g_bit[30].g_word[21].r_bit.Q ;
  wire \g_bit[30].g_word[22].r_bit.Q ;
  wire \g_bit[30].g_word[23].r_bit.Q ;
  wire \g_bit[30].g_word[24].r_bit.Q ;
  wire \g_bit[30].g_word[25].r_bit.Q ;
  wire \g_bit[30].g_word[26].r_bit.Q ;
  wire \g_bit[30].g_word[27].r_bit.Q ;
  wire \g_bit[30].g_word[28].r_bit.Q ;
  wire \g_bit[30].g_word[29].r_bit.Q ;
  wire \g_bit[30].g_word[2].r_bit.Q ;
  wire \g_bit[30].g_word[30].r_bit.Q ;
  wire \g_bit[30].g_word[31].r_bit.Q ;
  wire \g_bit[30].g_word[3].r_bit.Q ;
  wire \g_bit[30].g_word[4].r_bit.Q ;
  wire \g_bit[30].g_word[5].r_bit.Q ;
  wire \g_bit[30].g_word[6].r_bit.Q ;
  wire \g_bit[30].g_word[7].r_bit.Q ;
  wire \g_bit[30].g_word[8].r_bit.Q ;
  wire \g_bit[30].g_word[9].r_bit.Q ;
  wire \g_bit[30].r_rs1.D ;
  wire \g_bit[30].r_rs1.Q ;
  wire \g_bit[30].r_rs2.D ;
  wire \g_bit[30].r_rs2.Q ;
  wire \g_bit[31].g_word[10].r_bit.Q ;
  wire \g_bit[31].g_word[11].r_bit.Q ;
  wire \g_bit[31].g_word[12].r_bit.Q ;
  wire \g_bit[31].g_word[13].r_bit.Q ;
  wire \g_bit[31].g_word[14].r_bit.Q ;
  wire \g_bit[31].g_word[15].r_bit.Q ;
  wire \g_bit[31].g_word[16].r_bit.Q ;
  wire \g_bit[31].g_word[17].r_bit.Q ;
  wire \g_bit[31].g_word[18].r_bit.Q ;
  wire \g_bit[31].g_word[19].r_bit.Q ;
  wire \g_bit[31].g_word[1].r_bit.Q ;
  wire \g_bit[31].g_word[20].r_bit.Q ;
  wire \g_bit[31].g_word[21].r_bit.Q ;
  wire \g_bit[31].g_word[22].r_bit.Q ;
  wire \g_bit[31].g_word[23].r_bit.Q ;
  wire \g_bit[31].g_word[24].r_bit.Q ;
  wire \g_bit[31].g_word[25].r_bit.Q ;
  wire \g_bit[31].g_word[26].r_bit.Q ;
  wire \g_bit[31].g_word[27].r_bit.Q ;
  wire \g_bit[31].g_word[28].r_bit.Q ;
  wire \g_bit[31].g_word[29].r_bit.Q ;
  wire \g_bit[31].g_word[2].r_bit.Q ;
  wire \g_bit[31].g_word[30].r_bit.Q ;
  wire \g_bit[31].g_word[31].r_bit.Q ;
  wire \g_bit[31].g_word[3].r_bit.Q ;
  wire \g_bit[31].g_word[4].r_bit.Q ;
  wire \g_bit[31].g_word[5].r_bit.Q ;
  wire \g_bit[31].g_word[6].r_bit.Q ;
  wire \g_bit[31].g_word[7].r_bit.Q ;
  wire \g_bit[31].g_word[8].r_bit.Q ;
  wire \g_bit[31].g_word[9].r_bit.Q ;
  wire \g_bit[31].r_rs1.D ;
  wire \g_bit[31].r_rs1.Q ;
  wire \g_bit[31].r_rs2.D ;
  wire \g_bit[31].r_rs2.Q ;
  wire \g_bit[3].g_word[10].r_bit.Q ;
  wire \g_bit[3].g_word[11].r_bit.Q ;
  wire \g_bit[3].g_word[12].r_bit.Q ;
  wire \g_bit[3].g_word[13].r_bit.Q ;
  wire \g_bit[3].g_word[14].r_bit.Q ;
  wire \g_bit[3].g_word[15].r_bit.Q ;
  wire \g_bit[3].g_word[16].r_bit.Q ;
  wire \g_bit[3].g_word[17].r_bit.Q ;
  wire \g_bit[3].g_word[18].r_bit.Q ;
  wire \g_bit[3].g_word[19].r_bit.Q ;
  wire \g_bit[3].g_word[1].r_bit.Q ;
  wire \g_bit[3].g_word[20].r_bit.Q ;
  wire \g_bit[3].g_word[21].r_bit.Q ;
  wire \g_bit[3].g_word[22].r_bit.Q ;
  wire \g_bit[3].g_word[23].r_bit.Q ;
  wire \g_bit[3].g_word[24].r_bit.Q ;
  wire \g_bit[3].g_word[25].r_bit.Q ;
  wire \g_bit[3].g_word[26].r_bit.Q ;
  wire \g_bit[3].g_word[27].r_bit.Q ;
  wire \g_bit[3].g_word[28].r_bit.Q ;
  wire \g_bit[3].g_word[29].r_bit.Q ;
  wire \g_bit[3].g_word[2].r_bit.Q ;
  wire \g_bit[3].g_word[30].r_bit.Q ;
  wire \g_bit[3].g_word[31].r_bit.Q ;
  wire \g_bit[3].g_word[3].r_bit.Q ;
  wire \g_bit[3].g_word[4].r_bit.Q ;
  wire \g_bit[3].g_word[5].r_bit.Q ;
  wire \g_bit[3].g_word[6].r_bit.Q ;
  wire \g_bit[3].g_word[7].r_bit.Q ;
  wire \g_bit[3].g_word[8].r_bit.Q ;
  wire \g_bit[3].g_word[9].r_bit.Q ;
  wire \g_bit[3].r_rs1.D ;
  wire \g_bit[3].r_rs1.Q ;
  wire \g_bit[3].r_rs2.D ;
  wire \g_bit[3].r_rs2.Q ;
  wire \g_bit[4].g_word[10].r_bit.Q ;
  wire \g_bit[4].g_word[11].r_bit.Q ;
  wire \g_bit[4].g_word[12].r_bit.Q ;
  wire \g_bit[4].g_word[13].r_bit.Q ;
  wire \g_bit[4].g_word[14].r_bit.Q ;
  wire \g_bit[4].g_word[15].r_bit.Q ;
  wire \g_bit[4].g_word[16].r_bit.Q ;
  wire \g_bit[4].g_word[17].r_bit.Q ;
  wire \g_bit[4].g_word[18].r_bit.Q ;
  wire \g_bit[4].g_word[19].r_bit.Q ;
  wire \g_bit[4].g_word[1].r_bit.Q ;
  wire \g_bit[4].g_word[20].r_bit.Q ;
  wire \g_bit[4].g_word[21].r_bit.Q ;
  wire \g_bit[4].g_word[22].r_bit.Q ;
  wire \g_bit[4].g_word[23].r_bit.Q ;
  wire \g_bit[4].g_word[24].r_bit.Q ;
  wire \g_bit[4].g_word[25].r_bit.Q ;
  wire \g_bit[4].g_word[26].r_bit.Q ;
  wire \g_bit[4].g_word[27].r_bit.Q ;
  wire \g_bit[4].g_word[28].r_bit.Q ;
  wire \g_bit[4].g_word[29].r_bit.Q ;
  wire \g_bit[4].g_word[2].r_bit.Q ;
  wire \g_bit[4].g_word[30].r_bit.Q ;
  wire \g_bit[4].g_word[31].r_bit.Q ;
  wire \g_bit[4].g_word[3].r_bit.Q ;
  wire \g_bit[4].g_word[4].r_bit.Q ;
  wire \g_bit[4].g_word[5].r_bit.Q ;
  wire \g_bit[4].g_word[6].r_bit.Q ;
  wire \g_bit[4].g_word[7].r_bit.Q ;
  wire \g_bit[4].g_word[8].r_bit.Q ;
  wire \g_bit[4].g_word[9].r_bit.Q ;
  wire \g_bit[4].r_rs1.D ;
  wire \g_bit[4].r_rs1.Q ;
  wire \g_bit[4].r_rs2.D ;
  wire \g_bit[4].r_rs2.Q ;
  wire \g_bit[5].g_word[10].r_bit.Q ;
  wire \g_bit[5].g_word[11].r_bit.Q ;
  wire \g_bit[5].g_word[12].r_bit.Q ;
  wire \g_bit[5].g_word[13].r_bit.Q ;
  wire \g_bit[5].g_word[14].r_bit.Q ;
  wire \g_bit[5].g_word[15].r_bit.Q ;
  wire \g_bit[5].g_word[16].r_bit.Q ;
  wire \g_bit[5].g_word[17].r_bit.Q ;
  wire \g_bit[5].g_word[18].r_bit.Q ;
  wire \g_bit[5].g_word[19].r_bit.Q ;
  wire \g_bit[5].g_word[1].r_bit.Q ;
  wire \g_bit[5].g_word[20].r_bit.Q ;
  wire \g_bit[5].g_word[21].r_bit.Q ;
  wire \g_bit[5].g_word[22].r_bit.Q ;
  wire \g_bit[5].g_word[23].r_bit.Q ;
  wire \g_bit[5].g_word[24].r_bit.Q ;
  wire \g_bit[5].g_word[25].r_bit.Q ;
  wire \g_bit[5].g_word[26].r_bit.Q ;
  wire \g_bit[5].g_word[27].r_bit.Q ;
  wire \g_bit[5].g_word[28].r_bit.Q ;
  wire \g_bit[5].g_word[29].r_bit.Q ;
  wire \g_bit[5].g_word[2].r_bit.Q ;
  wire \g_bit[5].g_word[30].r_bit.Q ;
  wire \g_bit[5].g_word[31].r_bit.Q ;
  wire \g_bit[5].g_word[3].r_bit.Q ;
  wire \g_bit[5].g_word[4].r_bit.Q ;
  wire \g_bit[5].g_word[5].r_bit.Q ;
  wire \g_bit[5].g_word[6].r_bit.Q ;
  wire \g_bit[5].g_word[7].r_bit.Q ;
  wire \g_bit[5].g_word[8].r_bit.Q ;
  wire \g_bit[5].g_word[9].r_bit.Q ;
  wire \g_bit[5].r_rs1.D ;
  wire \g_bit[5].r_rs1.Q ;
  wire \g_bit[5].r_rs2.D ;
  wire \g_bit[5].r_rs2.Q ;
  wire \g_bit[6].g_word[10].r_bit.Q ;
  wire \g_bit[6].g_word[11].r_bit.Q ;
  wire \g_bit[6].g_word[12].r_bit.Q ;
  wire \g_bit[6].g_word[13].r_bit.Q ;
  wire \g_bit[6].g_word[14].r_bit.Q ;
  wire \g_bit[6].g_word[15].r_bit.Q ;
  wire \g_bit[6].g_word[16].r_bit.Q ;
  wire \g_bit[6].g_word[17].r_bit.Q ;
  wire \g_bit[6].g_word[18].r_bit.Q ;
  wire \g_bit[6].g_word[19].r_bit.Q ;
  wire \g_bit[6].g_word[1].r_bit.Q ;
  wire \g_bit[6].g_word[20].r_bit.Q ;
  wire \g_bit[6].g_word[21].r_bit.Q ;
  wire \g_bit[6].g_word[22].r_bit.Q ;
  wire \g_bit[6].g_word[23].r_bit.Q ;
  wire \g_bit[6].g_word[24].r_bit.Q ;
  wire \g_bit[6].g_word[25].r_bit.Q ;
  wire \g_bit[6].g_word[26].r_bit.Q ;
  wire \g_bit[6].g_word[27].r_bit.Q ;
  wire \g_bit[6].g_word[28].r_bit.Q ;
  wire \g_bit[6].g_word[29].r_bit.Q ;
  wire \g_bit[6].g_word[2].r_bit.Q ;
  wire \g_bit[6].g_word[30].r_bit.Q ;
  wire \g_bit[6].g_word[31].r_bit.Q ;
  wire \g_bit[6].g_word[3].r_bit.Q ;
  wire \g_bit[6].g_word[4].r_bit.Q ;
  wire \g_bit[6].g_word[5].r_bit.Q ;
  wire \g_bit[6].g_word[6].r_bit.Q ;
  wire \g_bit[6].g_word[7].r_bit.Q ;
  wire \g_bit[6].g_word[8].r_bit.Q ;
  wire \g_bit[6].g_word[9].r_bit.Q ;
  wire \g_bit[6].r_rs1.D ;
  wire \g_bit[6].r_rs1.Q ;
  wire \g_bit[6].r_rs2.D ;
  wire \g_bit[6].r_rs2.Q ;
  wire \g_bit[7].g_word[10].r_bit.Q ;
  wire \g_bit[7].g_word[11].r_bit.Q ;
  wire \g_bit[7].g_word[12].r_bit.Q ;
  wire \g_bit[7].g_word[13].r_bit.Q ;
  wire \g_bit[7].g_word[14].r_bit.Q ;
  wire \g_bit[7].g_word[15].r_bit.Q ;
  wire \g_bit[7].g_word[16].r_bit.Q ;
  wire \g_bit[7].g_word[17].r_bit.Q ;
  wire \g_bit[7].g_word[18].r_bit.Q ;
  wire \g_bit[7].g_word[19].r_bit.Q ;
  wire \g_bit[7].g_word[1].r_bit.Q ;
  wire \g_bit[7].g_word[20].r_bit.Q ;
  wire \g_bit[7].g_word[21].r_bit.Q ;
  wire \g_bit[7].g_word[22].r_bit.Q ;
  wire \g_bit[7].g_word[23].r_bit.Q ;
  wire \g_bit[7].g_word[24].r_bit.Q ;
  wire \g_bit[7].g_word[25].r_bit.Q ;
  wire \g_bit[7].g_word[26].r_bit.Q ;
  wire \g_bit[7].g_word[27].r_bit.Q ;
  wire \g_bit[7].g_word[28].r_bit.Q ;
  wire \g_bit[7].g_word[29].r_bit.Q ;
  wire \g_bit[7].g_word[2].r_bit.Q ;
  wire \g_bit[7].g_word[30].r_bit.Q ;
  wire \g_bit[7].g_word[31].r_bit.Q ;
  wire \g_bit[7].g_word[3].r_bit.Q ;
  wire \g_bit[7].g_word[4].r_bit.Q ;
  wire \g_bit[7].g_word[5].r_bit.Q ;
  wire \g_bit[7].g_word[6].r_bit.Q ;
  wire \g_bit[7].g_word[7].r_bit.Q ;
  wire \g_bit[7].g_word[8].r_bit.Q ;
  wire \g_bit[7].g_word[9].r_bit.Q ;
  wire \g_bit[7].r_rs1.D ;
  wire \g_bit[7].r_rs1.Q ;
  wire \g_bit[7].r_rs2.D ;
  wire \g_bit[7].r_rs2.Q ;
  wire \g_bit[8].g_word[10].r_bit.Q ;
  wire \g_bit[8].g_word[11].r_bit.Q ;
  wire \g_bit[8].g_word[12].r_bit.Q ;
  wire \g_bit[8].g_word[13].r_bit.Q ;
  wire \g_bit[8].g_word[14].r_bit.Q ;
  wire \g_bit[8].g_word[15].r_bit.Q ;
  wire \g_bit[8].g_word[16].r_bit.Q ;
  wire \g_bit[8].g_word[17].r_bit.Q ;
  wire \g_bit[8].g_word[18].r_bit.Q ;
  wire \g_bit[8].g_word[19].r_bit.Q ;
  wire \g_bit[8].g_word[1].r_bit.Q ;
  wire \g_bit[8].g_word[20].r_bit.Q ;
  wire \g_bit[8].g_word[21].r_bit.Q ;
  wire \g_bit[8].g_word[22].r_bit.Q ;
  wire \g_bit[8].g_word[23].r_bit.Q ;
  wire \g_bit[8].g_word[24].r_bit.Q ;
  wire \g_bit[8].g_word[25].r_bit.Q ;
  wire \g_bit[8].g_word[26].r_bit.Q ;
  wire \g_bit[8].g_word[27].r_bit.Q ;
  wire \g_bit[8].g_word[28].r_bit.Q ;
  wire \g_bit[8].g_word[29].r_bit.Q ;
  wire \g_bit[8].g_word[2].r_bit.Q ;
  wire \g_bit[8].g_word[30].r_bit.Q ;
  wire \g_bit[8].g_word[31].r_bit.Q ;
  wire \g_bit[8].g_word[3].r_bit.Q ;
  wire \g_bit[8].g_word[4].r_bit.Q ;
  wire \g_bit[8].g_word[5].r_bit.Q ;
  wire \g_bit[8].g_word[6].r_bit.Q ;
  wire \g_bit[8].g_word[7].r_bit.Q ;
  wire \g_bit[8].g_word[8].r_bit.Q ;
  wire \g_bit[8].g_word[9].r_bit.Q ;
  wire \g_bit[8].r_rs1.D ;
  wire \g_bit[8].r_rs1.Q ;
  wire \g_bit[8].r_rs2.D ;
  wire \g_bit[8].r_rs2.Q ;
  wire \g_bit[9].g_word[10].r_bit.Q ;
  wire \g_bit[9].g_word[11].r_bit.Q ;
  wire \g_bit[9].g_word[12].r_bit.Q ;
  wire \g_bit[9].g_word[13].r_bit.Q ;
  wire \g_bit[9].g_word[14].r_bit.Q ;
  wire \g_bit[9].g_word[15].r_bit.Q ;
  wire \g_bit[9].g_word[16].r_bit.Q ;
  wire \g_bit[9].g_word[17].r_bit.Q ;
  wire \g_bit[9].g_word[18].r_bit.Q ;
  wire \g_bit[9].g_word[19].r_bit.Q ;
  wire \g_bit[9].g_word[1].r_bit.Q ;
  wire \g_bit[9].g_word[20].r_bit.Q ;
  wire \g_bit[9].g_word[21].r_bit.Q ;
  wire \g_bit[9].g_word[22].r_bit.Q ;
  wire \g_bit[9].g_word[23].r_bit.Q ;
  wire \g_bit[9].g_word[24].r_bit.Q ;
  wire \g_bit[9].g_word[25].r_bit.Q ;
  wire \g_bit[9].g_word[26].r_bit.Q ;
  wire \g_bit[9].g_word[27].r_bit.Q ;
  wire \g_bit[9].g_word[28].r_bit.Q ;
  wire \g_bit[9].g_word[29].r_bit.Q ;
  wire \g_bit[9].g_word[2].r_bit.Q ;
  wire \g_bit[9].g_word[30].r_bit.Q ;
  wire \g_bit[9].g_word[31].r_bit.Q ;
  wire \g_bit[9].g_word[3].r_bit.Q ;
  wire \g_bit[9].g_word[4].r_bit.Q ;
  wire \g_bit[9].g_word[5].r_bit.Q ;
  wire \g_bit[9].g_word[6].r_bit.Q ;
  wire \g_bit[9].g_word[7].r_bit.Q ;
  wire \g_bit[9].g_word[8].r_bit.Q ;
  wire \g_bit[9].g_word[9].r_bit.Q ;
  wire \g_bit[9].r_rs1.D ;
  wire \g_bit[9].r_rs1.Q ;
  wire \g_bit[9].r_rs2.D ;
  wire \g_bit[9].r_rs2.Q ;
  input i_clk;
  wire i_clk;
  input [31:0] i_data;
  wire [31:0] i_data;
  input [4:0] i_rd;
  wire [4:0] i_rd;
  input i_reset_n;
  wire i_reset_n;
  input [4:0] i_rs1;
  wire [4:0] i_rs1;
  input [4:0] i_rs2;
  wire [4:0] i_rs2;
  input i_rs_valid;
  wire i_rs_valid;
  input i_write;
  wire i_write;
  output [31:0] o_data1;
  wire [31:0] o_data1;
  output [31:0] o_data2;
  wire [31:0] o_data2;
  wire \r_rs1[0].Q ;
  wire \r_rs1[1].Q ;
  wire \r_rs1[2].Q ;
  wire \r_rs1[3].Q ;
  wire \r_rs1[4].Q ;
  wire \r_rs2[0].Q ;
  wire \r_rs2[1].Q ;
  wire \r_rs2[2].Q ;
  wire \r_rs2[3].Q ;
  wire \r_rs2[4].Q ;
  wire[31:0] rs1;
  wire[31:0] rs2;
  sky130_fd_sc_hd__or2b_2 _2302_ (
    .A(rs1[3]),
    .B_N(rs1[2]),
    .X(_0002_)
  );
  sky130_fd_sc_hd__buf_1 _2303_ (
    .A(_0002_),
    .X(_0003_)
  );
  sky130_fd_sc_hd__buf_1 _2304_ (
    .A(_0003_),
    .X(_0004_)
  );
  sky130_fd_sc_hd__buf_1 _2306_ (
    .A(rs1[4]),
    .X(_0006_)
  );
  sky130_fd_sc_hd__buf_1 _2308_ (
    .A(rs1[1]),
    .X(_0008_)
  );
  sky130_fd_sc_hd__buf_1 _2310_ (
    .A(rs1[0]),
    .X(_0010_)
  );
  sky130_fd_sc_hd__or3_2 _2311_ (
    .A(_0006_),
    .B(_0008_),
    .C(_0010_),
    .X(_0011_)
  );
  sky130_fd_sc_hd__buf_1 _2312_ (
    .A(_0011_),
    .X(_0012_)
  );
  sky130_fd_sc_hd__nor2_2 _2313_ (
    .A(_0004_),
    .B(_0012_),
    .Y(_0013_)
  );
  sky130_fd_sc_hd__buf_1 _2314_ (
    .A(_0013_),
    .X(_0014_)
  );
  sky130_fd_sc_hd__nand2b_2 _2315_ (
    .A_N(rs1[2]),
    .B(rs1[3]),
    .Y(_0015_)
  );
  sky130_fd_sc_hd__buf_1 _2316_ (
    .A(_0015_),
    .X(_0016_)
  );
  sky130_fd_sc_hd__buf_1 _2317_ (
    .A(_0016_),
    .X(_0017_)
  );
  sky130_fd_sc_hd__nand3b_2 _2318_ (
    .A_N(_0010_),
    .B(_0008_),
    .C(_0006_),
    .Y(_0018_)
  );
  sky130_fd_sc_hd__buf_1 _2319_ (
    .A(_0018_),
    .X(_0019_)
  );
  sky130_fd_sc_hd__nor2_2 _2320_ (
    .A(_0017_),
    .B(_0019_),
    .Y(_0020_)
  );
  sky130_fd_sc_hd__buf_1 _2321_ (
    .A(_0020_),
    .X(_0021_)
  );
  sky130_fd_sc_hd__and2_2 _2322_ (
    .A(rs1[3]),
    .B(rs1[2]),
    .X(_0022_)
  );
  sky130_fd_sc_hd__buf_1 _2323_ (
    .A(_0022_),
    .X(_0023_)
  );
  sky130_fd_sc_hd__and3b_2 _2324_ (
    .A_N(_0010_),
    .B(_0008_),
    .C(_0006_),
    .X(_0024_)
  );
  sky130_fd_sc_hd__buf_1 _2325_ (
    .A(_0024_),
    .X(_0025_)
  );
  sky130_fd_sc_hd__or3b_2 _2326_ (
    .A(_0008_),
    .B(_0010_),
    .C_N(_0006_),
    .X(_0026_)
  );
  sky130_fd_sc_hd__nand2_2 _2327_ (
    .A(rs1[3]),
    .B(rs1[2]),
    .Y(_0027_)
  );
  sky130_fd_sc_hd__buf_1 _2328_ (
    .A(_0027_),
    .X(_0028_)
  );
  sky130_fd_sc_hd__nor2_2 _2329_ (
    .A(_0026_),
    .B(_0028_),
    .Y(_0029_)
  );
  sky130_fd_sc_hd__buf_1 _2330_ (
    .A(_0029_),
    .X(_0030_)
  );
  sky130_fd_sc_hd__a32o_2 _2331_ (
    .A1(\g_bit[31].g_word[30].r_bit.Q ),
    .A2(_0023_),
    .A3(_0025_),
    .B1(_0030_),
    .B2(\g_bit[31].g_word[28].r_bit.Q ),
    .X(_0031_)
  );
  sky130_fd_sc_hd__a221o_2 _2332_ (
    .A1(\g_bit[31].g_word[4].r_bit.Q ),
    .A2(_0014_),
    .B1(_0021_),
    .B2(\g_bit[31].g_word[26].r_bit.Q ),
    .C1(_0031_),
    .X(_0032_)
  );
  sky130_fd_sc_hd__nand3b_2 _2333_ (
    .A_N(_0008_),
    .B(_0010_),
    .C(_0006_),
    .Y(_0033_)
  );
  sky130_fd_sc_hd__nor2_2 _2334_ (
    .A(_0017_),
    .B(_0033_),
    .Y(_0034_)
  );
  sky130_fd_sc_hd__buf_1 _2335_ (
    .A(_0034_),
    .X(_0035_)
  );
  sky130_fd_sc_hd__nand3_2 _2336_ (
    .A(_0006_),
    .B(_0008_),
    .C(_0010_),
    .Y(_0036_)
  );
  sky130_fd_sc_hd__buf_1 _2337_ (
    .A(_0028_),
    .X(_0037_)
  );
  sky130_fd_sc_hd__nor2_2 _2338_ (
    .A(_0036_),
    .B(_0037_),
    .Y(_0038_)
  );
  sky130_fd_sc_hd__buf_1 _2339_ (
    .A(_0038_),
    .X(_0039_)
  );
  sky130_fd_sc_hd__or3b_2 _2340_ (
    .A(_0006_),
    .B(_0008_),
    .C_N(_0010_),
    .X(_0040_)
  );
  sky130_fd_sc_hd__buf_1 _2341_ (
    .A(_0040_),
    .X(_0041_)
  );
  sky130_fd_sc_hd__nor2_2 _2342_ (
    .A(_0003_),
    .B(_0041_),
    .Y(_0042_)
  );
  sky130_fd_sc_hd__buf_1 _2343_ (
    .A(_0042_),
    .X(_0043_)
  );
  sky130_fd_sc_hd__or2_2 _2344_ (
    .A(rs1[3]),
    .B(rs1[2]),
    .X(_0044_)
  );
  sky130_fd_sc_hd__buf_1 _2345_ (
    .A(_0044_),
    .X(_0045_)
  );
  sky130_fd_sc_hd__buf_1 _2346_ (
    .A(_0045_),
    .X(_0046_)
  );
  sky130_fd_sc_hd__or3b_2 _2347_ (
    .A(rs1[4]),
    .B(rs1[0]),
    .C_N(rs1[1]),
    .X(_0047_)
  );
  sky130_fd_sc_hd__buf_1 _2348_ (
    .A(_0047_),
    .X(_0048_)
  );
  sky130_fd_sc_hd__nor2_2 _2349_ (
    .A(_0046_),
    .B(_0048_),
    .Y(_0049_)
  );
  sky130_fd_sc_hd__buf_1 _2350_ (
    .A(_0049_),
    .X(_0050_)
  );
  sky130_fd_sc_hd__a22o_2 _2351_ (
    .A1(\g_bit[31].g_word[5].r_bit.Q ),
    .A2(_0043_),
    .B1(_0050_),
    .B2(\g_bit[31].g_word[2].r_bit.Q ),
    .X(_0051_)
  );
  sky130_fd_sc_hd__a221o_2 _2352_ (
    .A1(\g_bit[31].g_word[25].r_bit.Q ),
    .A2(_0035_),
    .B1(_0039_),
    .B2(\g_bit[31].g_word[31].r_bit.Q ),
    .C1(_0051_),
    .X(_0052_)
  );
  sky130_fd_sc_hd__nor2_2 _2353_ (
    .A(_0028_),
    .B(_0041_),
    .Y(_0053_)
  );
  sky130_fd_sc_hd__buf_1 _2354_ (
    .A(_0053_),
    .X(_0054_)
  );
  sky130_fd_sc_hd__nand3b_2 _2355_ (
    .A_N(_0006_),
    .B(_0008_),
    .C(_0010_),
    .Y(_0055_)
  );
  sky130_fd_sc_hd__nor2_2 _2356_ (
    .A(_0055_),
    .B(_0028_),
    .Y(_0056_)
  );
  sky130_fd_sc_hd__buf_1 _2357_ (
    .A(_0056_),
    .X(_0057_)
  );
  sky130_fd_sc_hd__a22o_2 _2358_ (
    .A1(\g_bit[31].g_word[13].r_bit.Q ),
    .A2(_0054_),
    .B1(_0057_),
    .B2(\g_bit[31].g_word[15].r_bit.Q ),
    .X(_0058_)
  );
  sky130_fd_sc_hd__nor2_2 _2359_ (
    .A(_0015_),
    .B(_0055_),
    .Y(_0059_)
  );
  sky130_fd_sc_hd__buf_1 _2360_ (
    .A(_0059_),
    .X(_0060_)
  );
  sky130_fd_sc_hd__nor2_2 _2361_ (
    .A(_0026_),
    .B(_0003_),
    .Y(_0061_)
  );
  sky130_fd_sc_hd__buf_1 _2362_ (
    .A(_0061_),
    .X(_0062_)
  );
  sky130_fd_sc_hd__a22o_2 _2363_ (
    .A1(\g_bit[31].g_word[11].r_bit.Q ),
    .A2(_0060_),
    .B1(_0062_),
    .B2(\g_bit[31].g_word[20].r_bit.Q ),
    .X(_0063_)
  );
  sky130_fd_sc_hd__nor2_2 _2364_ (
    .A(_0036_),
    .B(_0045_),
    .Y(_0064_)
  );
  sky130_fd_sc_hd__buf_1 _2365_ (
    .A(_0064_),
    .X(_0065_)
  );
  sky130_fd_sc_hd__nor2_2 _2366_ (
    .A(_0033_),
    .B(_0003_),
    .Y(_0066_)
  );
  sky130_fd_sc_hd__buf_1 _2367_ (
    .A(_0066_),
    .X(_0067_)
  );
  sky130_fd_sc_hd__a22o_2 _2368_ (
    .A1(\g_bit[31].g_word[19].r_bit.Q ),
    .A2(_0065_),
    .B1(_0067_),
    .B2(\g_bit[31].g_word[21].r_bit.Q ),
    .X(_0068_)
  );
  sky130_fd_sc_hd__nor2_2 _2369_ (
    .A(_0045_),
    .B(_0033_),
    .Y(_0069_)
  );
  sky130_fd_sc_hd__buf_1 _2370_ (
    .A(_0069_),
    .X(_0070_)
  );
  sky130_fd_sc_hd__nor2_2 _2371_ (
    .A(_0028_),
    .B(_0011_),
    .Y(_0071_)
  );
  sky130_fd_sc_hd__buf_1 _2372_ (
    .A(_0071_),
    .X(_0072_)
  );
  sky130_fd_sc_hd__a22o_2 _2373_ (
    .A1(\g_bit[31].g_word[17].r_bit.Q ),
    .A2(_0070_),
    .B1(_0072_),
    .B2(\g_bit[31].g_word[12].r_bit.Q ),
    .X(_0073_)
  );
  sky130_fd_sc_hd__or4_2 _2374_ (
    .A(_0058_),
    .B(_0063_),
    .C(_0068_),
    .D(_0073_),
    .X(_0074_)
  );
  sky130_fd_sc_hd__nor2_2 _2375_ (
    .A(_0033_),
    .B(_0027_),
    .Y(_0075_)
  );
  sky130_fd_sc_hd__buf_1 _2376_ (
    .A(_0075_),
    .X(_0076_)
  );
  sky130_fd_sc_hd__nor2b_2 _2377_ (
    .A(rs1[2]),
    .B_N(rs1[3]),
    .Y(_0077_)
  );
  sky130_fd_sc_hd__nor3b_2 _2378_ (
    .A(_0008_),
    .B(_0010_),
    .C_N(_0006_),
    .Y(_0078_)
  );
  sky130_fd_sc_hd__and3_2 _2379_ (
    .A(\g_bit[31].g_word[24].r_bit.Q ),
    .B(_0077_),
    .C(_0078_),
    .X(_0079_)
  );
  sky130_fd_sc_hd__inv_2 _2380_ (
    .A(\g_bit[31].g_word[7].r_bit.Q ),
    .Y(_0080_)
  );
  sky130_fd_sc_hd__buf_1 _2381_ (
    .A(_0055_),
    .X(_0081_)
  );
  sky130_fd_sc_hd__buf_1 _2382_ (
    .A(_0081_),
    .X(_0082_)
  );
  sky130_fd_sc_hd__nor3_2 _2383_ (
    .A(_0080_),
    .B(_0082_),
    .C(_0004_),
    .Y(_0083_)
  );
  sky130_fd_sc_hd__inv_2 _2384_ (
    .A(\g_bit[31].g_word[3].r_bit.Q ),
    .Y(_0084_)
  );
  sky130_fd_sc_hd__buf_1 _2385_ (
    .A(_0045_),
    .X(_0085_)
  );
  sky130_fd_sc_hd__buf_1 _2386_ (
    .A(_0081_),
    .X(_0086_)
  );
  sky130_fd_sc_hd__nor3_2 _2387_ (
    .A(_0084_),
    .B(_0085_),
    .C(_0086_),
    .Y(_0087_)
  );
  sky130_fd_sc_hd__a2111o_2 _2388_ (
    .A1(\g_bit[31].g_word[29].r_bit.Q ),
    .A2(_0076_),
    .B1(_0079_),
    .C1(_0083_),
    .D1(_0087_),
    .X(_0088_)
  );
  sky130_fd_sc_hd__nor2_2 _2389_ (
    .A(_0003_),
    .B(_0047_),
    .Y(_0089_)
  );
  sky130_fd_sc_hd__buf_1 _2390_ (
    .A(_0089_),
    .X(_0090_)
  );
  sky130_fd_sc_hd__nor2_2 _2391_ (
    .A(_0045_),
    .B(_0041_),
    .Y(_0091_)
  );
  sky130_fd_sc_hd__buf_1 _2392_ (
    .A(_0091_),
    .X(_0092_)
  );
  sky130_fd_sc_hd__and3_2 _2393_ (
    .A(_0006_),
    .B(_0008_),
    .C(_0010_),
    .X(_0093_)
  );
  sky130_fd_sc_hd__buf_1 _2394_ (
    .A(_0093_),
    .X(_0094_)
  );
  sky130_fd_sc_hd__buf_1 _2395_ (
    .A(_0077_),
    .X(_0095_)
  );
  sky130_fd_sc_hd__and3_2 _2396_ (
    .A(\g_bit[31].g_word[27].r_bit.Q ),
    .B(_0094_),
    .C(_0095_),
    .X(_0096_)
  );
  sky130_fd_sc_hd__a221o_2 _2397_ (
    .A1(\g_bit[31].g_word[6].r_bit.Q ),
    .A2(_0090_),
    .B1(_0092_),
    .B2(\g_bit[31].g_word[1].r_bit.Q ),
    .C1(_0096_),
    .X(_0097_)
  );
  sky130_fd_sc_hd__inv_2 _2398_ (
    .A(\g_bit[31].g_word[23].r_bit.Q ),
    .Y(_0098_)
  );
  sky130_fd_sc_hd__or2_2 _2399_ (
    .A(_0036_),
    .B(_0002_),
    .X(_0099_)
  );
  sky130_fd_sc_hd__buf_1 _2400_ (
    .A(_0099_),
    .X(_0100_)
  );
  sky130_fd_sc_hd__buf_1 _2401_ (
    .A(_0100_),
    .X(_0101_)
  );
  sky130_fd_sc_hd__inv_2 _2402_ (
    .A(\g_bit[31].g_word[8].r_bit.Q ),
    .Y(_0102_)
  );
  sky130_fd_sc_hd__buf_1 _2403_ (
    .A(_0015_),
    .X(_0103_)
  );
  sky130_fd_sc_hd__or3_2 _2404_ (
    .A(_0102_),
    .B(_0103_),
    .C(_0011_),
    .X(_0104_)
  );
  sky130_fd_sc_hd__inv_2 _2405_ (
    .A(\g_bit[31].g_word[10].r_bit.Q ),
    .Y(_0105_)
  );
  sky130_fd_sc_hd__buf_1 _2406_ (
    .A(_0015_),
    .X(_0106_)
  );
  sky130_fd_sc_hd__buf_1 _2407_ (
    .A(_0047_),
    .X(_0107_)
  );
  sky130_fd_sc_hd__or3_2 _2408_ (
    .A(_0105_),
    .B(_0106_),
    .C(_0107_),
    .X(_0108_)
  );
  sky130_fd_sc_hd__inv_2 _2409_ (
    .A(\g_bit[31].g_word[9].r_bit.Q ),
    .Y(_0109_)
  );
  sky130_fd_sc_hd__buf_1 _2410_ (
    .A(_0041_),
    .X(_0110_)
  );
  sky130_fd_sc_hd__or3_2 _2411_ (
    .A(_0109_),
    .B(_0017_),
    .C(_0110_),
    .X(_0111_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2412_ (
    .A1(_0098_),
    .A2(_0101_),
    .B1(_0104_),
    .C1(_0108_),
    .D1(_0111_),
    .Y(_0112_)
  );
  sky130_fd_sc_hd__inv_2 _2413_ (
    .A(\g_bit[31].g_word[22].r_bit.Q ),
    .Y(_0113_)
  );
  sky130_fd_sc_hd__or2_2 _2414_ (
    .A(_0002_),
    .B(_0018_),
    .X(_0114_)
  );
  sky130_fd_sc_hd__buf_1 _2415_ (
    .A(_0114_),
    .X(_0115_)
  );
  sky130_fd_sc_hd__buf_1 _2416_ (
    .A(_0115_),
    .X(_0116_)
  );
  sky130_fd_sc_hd__inv_2 _2417_ (
    .A(\g_bit[31].g_word[18].r_bit.Q ),
    .Y(_0117_)
  );
  sky130_fd_sc_hd__buf_1 _2418_ (
    .A(_0045_),
    .X(_0118_)
  );
  sky130_fd_sc_hd__or3_2 _2419_ (
    .A(_0117_),
    .B(_0118_),
    .C(_0018_),
    .X(_0119_)
  );
  sky130_fd_sc_hd__inv_2 _2420_ (
    .A(\g_bit[31].g_word[16].r_bit.Q ),
    .Y(_0120_)
  );
  sky130_fd_sc_hd__buf_1 _2421_ (
    .A(_0026_),
    .X(_0121_)
  );
  sky130_fd_sc_hd__or3_2 _2422_ (
    .A(_0120_),
    .B(_0118_),
    .C(_0121_),
    .X(_0122_)
  );
  sky130_fd_sc_hd__inv_2 _2423_ (
    .A(\g_bit[31].g_word[14].r_bit.Q ),
    .Y(_0123_)
  );
  sky130_fd_sc_hd__buf_1 _2424_ (
    .A(_0048_),
    .X(_0124_)
  );
  sky130_fd_sc_hd__or3_2 _2425_ (
    .A(_0123_),
    .B(_0124_),
    .C(_0037_),
    .X(_0125_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2426_ (
    .A1(_0113_),
    .A2(_0116_),
    .B1(_0119_),
    .C1(_0122_),
    .D1(_0125_),
    .Y(_0126_)
  );
  sky130_fd_sc_hd__or4_2 _2427_ (
    .A(_0088_),
    .B(_0097_),
    .C(_0112_),
    .D(_0126_),
    .X(_0127_)
  );
  sky130_fd_sc_hd__or4_2 _2428_ (
    .A(_0032_),
    .B(_0052_),
    .C(_0074_),
    .D(_0127_),
    .X(_0128_)
  );
  sky130_fd_sc_hd__buf_1 _2429_ (
    .A(_0128_),
    .X(\g_bit[31].r_rs1.D )
  );
  sky130_fd_sc_hd__or2b_2 _2432_ (
    .A(rs2[3]),
    .B_N(rs2[2]),
    .X(_0131_)
  );
  sky130_fd_sc_hd__buf_1 _2433_ (
    .A(_0131_),
    .X(_0132_)
  );
  sky130_fd_sc_hd__buf_1 _2434_ (
    .A(_0132_),
    .X(_0133_)
  );
  sky130_fd_sc_hd__buf_1 _2436_ (
    .A(rs2[4]),
    .X(_0135_)
  );
  sky130_fd_sc_hd__buf_1 _2438_ (
    .A(rs2[1]),
    .X(_0137_)
  );
  sky130_fd_sc_hd__buf_1 _2440_ (
    .A(rs2[0]),
    .X(_0139_)
  );
  sky130_fd_sc_hd__or3_2 _2441_ (
    .A(_0135_),
    .B(_0137_),
    .C(_0139_),
    .X(_0140_)
  );
  sky130_fd_sc_hd__buf_1 _2442_ (
    .A(_0140_),
    .X(_0141_)
  );
  sky130_fd_sc_hd__nor2_2 _2443_ (
    .A(_0133_),
    .B(_0141_),
    .Y(_0142_)
  );
  sky130_fd_sc_hd__buf_1 _2444_ (
    .A(_0142_),
    .X(_0143_)
  );
  sky130_fd_sc_hd__nand2b_2 _2445_ (
    .A_N(rs2[2]),
    .B(_0129_),
    .Y(_0144_)
  );
  sky130_fd_sc_hd__buf_1 _2446_ (
    .A(_0144_),
    .X(_0145_)
  );
  sky130_fd_sc_hd__buf_1 _2447_ (
    .A(_0145_),
    .X(_0146_)
  );
  sky130_fd_sc_hd__nand3b_2 _2448_ (
    .A_N(_0139_),
    .B(_0137_),
    .C(_0135_),
    .Y(_0147_)
  );
  sky130_fd_sc_hd__buf_1 _2449_ (
    .A(_0147_),
    .X(_0148_)
  );
  sky130_fd_sc_hd__nor2_2 _2450_ (
    .A(_0146_),
    .B(_0148_),
    .Y(_0149_)
  );
  sky130_fd_sc_hd__buf_1 _2451_ (
    .A(_0149_),
    .X(_0150_)
  );
  sky130_fd_sc_hd__and2_2 _2452_ (
    .A(_0129_),
    .B(rs2[2]),
    .X(_0151_)
  );
  sky130_fd_sc_hd__buf_1 _2453_ (
    .A(_0151_),
    .X(_0152_)
  );
  sky130_fd_sc_hd__and3b_2 _2454_ (
    .A_N(_0139_),
    .B(_0137_),
    .C(_0135_),
    .X(_0153_)
  );
  sky130_fd_sc_hd__buf_1 _2455_ (
    .A(_0153_),
    .X(_0154_)
  );
  sky130_fd_sc_hd__or3b_2 _2456_ (
    .A(_0137_),
    .B(_0139_),
    .C_N(_0135_),
    .X(_0155_)
  );
  sky130_fd_sc_hd__nand2_2 _2457_ (
    .A(_0129_),
    .B(rs2[2]),
    .Y(_0156_)
  );
  sky130_fd_sc_hd__buf_1 _2458_ (
    .A(_0156_),
    .X(_0157_)
  );
  sky130_fd_sc_hd__nor2_2 _2459_ (
    .A(_0155_),
    .B(_0157_),
    .Y(_0158_)
  );
  sky130_fd_sc_hd__buf_1 _2460_ (
    .A(_0158_),
    .X(_0159_)
  );
  sky130_fd_sc_hd__a32o_2 _2461_ (
    .A1(\g_bit[31].g_word[30].r_bit.Q ),
    .A2(_0152_),
    .A3(_0154_),
    .B1(_0159_),
    .B2(\g_bit[31].g_word[28].r_bit.Q ),
    .X(_0160_)
  );
  sky130_fd_sc_hd__a221o_2 _2462_ (
    .A1(\g_bit[31].g_word[4].r_bit.Q ),
    .A2(_0143_),
    .B1(_0150_),
    .B2(\g_bit[31].g_word[26].r_bit.Q ),
    .C1(_0160_),
    .X(_0161_)
  );
  sky130_fd_sc_hd__nand3b_2 _2463_ (
    .A_N(_0137_),
    .B(_0139_),
    .C(_0135_),
    .Y(_0162_)
  );
  sky130_fd_sc_hd__nor2_2 _2464_ (
    .A(_0146_),
    .B(_0162_),
    .Y(_0163_)
  );
  sky130_fd_sc_hd__buf_1 _2465_ (
    .A(_0163_),
    .X(_0164_)
  );
  sky130_fd_sc_hd__nand3_2 _2466_ (
    .A(_0135_),
    .B(_0137_),
    .C(_0139_),
    .Y(_0165_)
  );
  sky130_fd_sc_hd__buf_1 _2467_ (
    .A(_0157_),
    .X(_0166_)
  );
  sky130_fd_sc_hd__nor2_2 _2468_ (
    .A(_0165_),
    .B(_0166_),
    .Y(_0167_)
  );
  sky130_fd_sc_hd__buf_1 _2469_ (
    .A(_0167_),
    .X(_0168_)
  );
  sky130_fd_sc_hd__or3b_2 _2470_ (
    .A(_0135_),
    .B(_0137_),
    .C_N(_0139_),
    .X(_0169_)
  );
  sky130_fd_sc_hd__buf_1 _2471_ (
    .A(_0169_),
    .X(_0170_)
  );
  sky130_fd_sc_hd__nor2_2 _2472_ (
    .A(_0132_),
    .B(_0170_),
    .Y(_0171_)
  );
  sky130_fd_sc_hd__buf_1 _2473_ (
    .A(_0171_),
    .X(_0172_)
  );
  sky130_fd_sc_hd__or2_2 _2474_ (
    .A(_0129_),
    .B(rs2[2]),
    .X(_0173_)
  );
  sky130_fd_sc_hd__buf_1 _2475_ (
    .A(_0173_),
    .X(_0174_)
  );
  sky130_fd_sc_hd__buf_1 _2476_ (
    .A(_0174_),
    .X(_0175_)
  );
  sky130_fd_sc_hd__or3b_2 _2477_ (
    .A(rs2[4]),
    .B(rs2[0]),
    .C_N(rs2[1]),
    .X(_0176_)
  );
  sky130_fd_sc_hd__buf_1 _2478_ (
    .A(_0176_),
    .X(_0177_)
  );
  sky130_fd_sc_hd__nor2_2 _2479_ (
    .A(_0175_),
    .B(_0177_),
    .Y(_0178_)
  );
  sky130_fd_sc_hd__buf_1 _2480_ (
    .A(_0178_),
    .X(_0179_)
  );
  sky130_fd_sc_hd__a22o_2 _2481_ (
    .A1(\g_bit[31].g_word[5].r_bit.Q ),
    .A2(_0172_),
    .B1(_0179_),
    .B2(\g_bit[31].g_word[2].r_bit.Q ),
    .X(_0180_)
  );
  sky130_fd_sc_hd__a221o_2 _2482_ (
    .A1(\g_bit[31].g_word[25].r_bit.Q ),
    .A2(_0164_),
    .B1(_0168_),
    .B2(\g_bit[31].g_word[31].r_bit.Q ),
    .C1(_0180_),
    .X(_0181_)
  );
  sky130_fd_sc_hd__nor2_2 _2483_ (
    .A(_0157_),
    .B(_0170_),
    .Y(_0182_)
  );
  sky130_fd_sc_hd__buf_1 _2484_ (
    .A(_0182_),
    .X(_0183_)
  );
  sky130_fd_sc_hd__nand3b_2 _2485_ (
    .A_N(_0135_),
    .B(_0137_),
    .C(_0139_),
    .Y(_0184_)
  );
  sky130_fd_sc_hd__nor2_2 _2486_ (
    .A(_0184_),
    .B(_0157_),
    .Y(_0185_)
  );
  sky130_fd_sc_hd__buf_1 _2487_ (
    .A(_0185_),
    .X(_0186_)
  );
  sky130_fd_sc_hd__a22o_2 _2488_ (
    .A1(\g_bit[31].g_word[13].r_bit.Q ),
    .A2(_0183_),
    .B1(_0186_),
    .B2(\g_bit[31].g_word[15].r_bit.Q ),
    .X(_0187_)
  );
  sky130_fd_sc_hd__nor2_2 _2489_ (
    .A(_0132_),
    .B(_0155_),
    .Y(_0188_)
  );
  sky130_fd_sc_hd__buf_1 _2490_ (
    .A(_0188_),
    .X(_0189_)
  );
  sky130_fd_sc_hd__nor2_2 _2491_ (
    .A(_0184_),
    .B(_0144_),
    .Y(_0190_)
  );
  sky130_fd_sc_hd__buf_1 _2492_ (
    .A(_0190_),
    .X(_0191_)
  );
  sky130_fd_sc_hd__a22o_2 _2493_ (
    .A1(\g_bit[31].g_word[20].r_bit.Q ),
    .A2(_0189_),
    .B1(_0191_),
    .B2(\g_bit[31].g_word[11].r_bit.Q ),
    .X(_0192_)
  );
  sky130_fd_sc_hd__nor2_2 _2494_ (
    .A(_0165_),
    .B(_0174_),
    .Y(_0193_)
  );
  sky130_fd_sc_hd__buf_1 _2495_ (
    .A(_0193_),
    .X(_0194_)
  );
  sky130_fd_sc_hd__nor2_2 _2496_ (
    .A(_0132_),
    .B(_0162_),
    .Y(_0195_)
  );
  sky130_fd_sc_hd__buf_1 _2497_ (
    .A(_0195_),
    .X(_0196_)
  );
  sky130_fd_sc_hd__a22o_2 _2498_ (
    .A1(\g_bit[31].g_word[19].r_bit.Q ),
    .A2(_0194_),
    .B1(_0196_),
    .B2(\g_bit[31].g_word[21].r_bit.Q ),
    .X(_0197_)
  );
  sky130_fd_sc_hd__nor2_2 _2499_ (
    .A(_0174_),
    .B(_0162_),
    .Y(_0198_)
  );
  sky130_fd_sc_hd__buf_1 _2500_ (
    .A(_0198_),
    .X(_0199_)
  );
  sky130_fd_sc_hd__nor2_2 _2501_ (
    .A(_0157_),
    .B(_0140_),
    .Y(_0200_)
  );
  sky130_fd_sc_hd__buf_1 _2502_ (
    .A(_0200_),
    .X(_0201_)
  );
  sky130_fd_sc_hd__a22o_2 _2503_ (
    .A1(\g_bit[31].g_word[17].r_bit.Q ),
    .A2(_0199_),
    .B1(_0201_),
    .B2(\g_bit[31].g_word[12].r_bit.Q ),
    .X(_0202_)
  );
  sky130_fd_sc_hd__or4_2 _2504_ (
    .A(_0187_),
    .B(_0192_),
    .C(_0197_),
    .D(_0202_),
    .X(_0203_)
  );
  sky130_fd_sc_hd__nor2_2 _2505_ (
    .A(_0156_),
    .B(_0162_),
    .Y(_0204_)
  );
  sky130_fd_sc_hd__buf_1 _2506_ (
    .A(_0204_),
    .X(_0205_)
  );
  sky130_fd_sc_hd__nor3b_2 _2507_ (
    .A(_0137_),
    .B(_0139_),
    .C_N(_0135_),
    .Y(_0206_)
  );
  sky130_fd_sc_hd__nor2b_2 _2508_ (
    .A(rs2[2]),
    .B_N(_0129_),
    .Y(_0207_)
  );
  sky130_fd_sc_hd__and3_2 _2509_ (
    .A(\g_bit[31].g_word[24].r_bit.Q ),
    .B(_0206_),
    .C(_0207_),
    .X(_0208_)
  );
  sky130_fd_sc_hd__buf_1 _2510_ (
    .A(_0184_),
    .X(_0209_)
  );
  sky130_fd_sc_hd__buf_1 _2511_ (
    .A(_0209_),
    .X(_0210_)
  );
  sky130_fd_sc_hd__nor3_2 _2512_ (
    .A(_0080_),
    .B(_0133_),
    .C(_0210_),
    .Y(_0211_)
  );
  sky130_fd_sc_hd__buf_1 _2513_ (
    .A(_0174_),
    .X(_0212_)
  );
  sky130_fd_sc_hd__nor3_2 _2514_ (
    .A(_0084_),
    .B(_0212_),
    .C(_0210_),
    .Y(_0213_)
  );
  sky130_fd_sc_hd__a2111o_2 _2515_ (
    .A1(\g_bit[31].g_word[29].r_bit.Q ),
    .A2(_0205_),
    .B1(_0208_),
    .C1(_0211_),
    .D1(_0213_),
    .X(_0214_)
  );
  sky130_fd_sc_hd__nor2_2 _2516_ (
    .A(_0132_),
    .B(_0176_),
    .Y(_0215_)
  );
  sky130_fd_sc_hd__buf_1 _2517_ (
    .A(_0215_),
    .X(_0216_)
  );
  sky130_fd_sc_hd__nor2_2 _2518_ (
    .A(_0174_),
    .B(_0170_),
    .Y(_0217_)
  );
  sky130_fd_sc_hd__buf_1 _2519_ (
    .A(_0217_),
    .X(_0218_)
  );
  sky130_fd_sc_hd__and3_2 _2520_ (
    .A(_0135_),
    .B(_0137_),
    .C(_0139_),
    .X(_0219_)
  );
  sky130_fd_sc_hd__buf_1 _2521_ (
    .A(_0219_),
    .X(_0220_)
  );
  sky130_fd_sc_hd__buf_1 _2522_ (
    .A(_0207_),
    .X(_0221_)
  );
  sky130_fd_sc_hd__and3_2 _2523_ (
    .A(\g_bit[31].g_word[27].r_bit.Q ),
    .B(_0220_),
    .C(_0221_),
    .X(_0222_)
  );
  sky130_fd_sc_hd__a221o_2 _2524_ (
    .A1(\g_bit[31].g_word[6].r_bit.Q ),
    .A2(_0216_),
    .B1(_0218_),
    .B2(\g_bit[31].g_word[1].r_bit.Q ),
    .C1(_0222_),
    .X(_0223_)
  );
  sky130_fd_sc_hd__or2_2 _2525_ (
    .A(_0131_),
    .B(_0165_),
    .X(_0224_)
  );
  sky130_fd_sc_hd__buf_1 _2526_ (
    .A(_0224_),
    .X(_0225_)
  );
  sky130_fd_sc_hd__buf_1 _2527_ (
    .A(_0225_),
    .X(_0226_)
  );
  sky130_fd_sc_hd__buf_1 _2528_ (
    .A(_0144_),
    .X(_0227_)
  );
  sky130_fd_sc_hd__or3_2 _2529_ (
    .A(_0102_),
    .B(_0227_),
    .C(_0140_),
    .X(_0228_)
  );
  sky130_fd_sc_hd__buf_1 _2530_ (
    .A(_0144_),
    .X(_0229_)
  );
  sky130_fd_sc_hd__buf_1 _2531_ (
    .A(_0176_),
    .X(_0230_)
  );
  sky130_fd_sc_hd__or3_2 _2532_ (
    .A(_0105_),
    .B(_0229_),
    .C(_0230_),
    .X(_0231_)
  );
  sky130_fd_sc_hd__buf_1 _2533_ (
    .A(_0170_),
    .X(_0232_)
  );
  sky130_fd_sc_hd__or3_2 _2534_ (
    .A(_0109_),
    .B(_0146_),
    .C(_0232_),
    .X(_0233_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2535_ (
    .A1(_0098_),
    .A2(_0226_),
    .B1(_0228_),
    .C1(_0231_),
    .D1(_0233_),
    .Y(_0234_)
  );
  sky130_fd_sc_hd__or2_2 _2536_ (
    .A(_0131_),
    .B(_0147_),
    .X(_0235_)
  );
  sky130_fd_sc_hd__buf_1 _2537_ (
    .A(_0235_),
    .X(_0236_)
  );
  sky130_fd_sc_hd__buf_1 _2538_ (
    .A(_0236_),
    .X(_0237_)
  );
  sky130_fd_sc_hd__or3_2 _2539_ (
    .A(_0117_),
    .B(_0175_),
    .C(_0147_),
    .X(_0238_)
  );
  sky130_fd_sc_hd__buf_1 _2540_ (
    .A(_0155_),
    .X(_0239_)
  );
  sky130_fd_sc_hd__buf_1 _2541_ (
    .A(_0174_),
    .X(_0240_)
  );
  sky130_fd_sc_hd__or3_2 _2542_ (
    .A(_0120_),
    .B(_0239_),
    .C(_0240_),
    .X(_0241_)
  );
  sky130_fd_sc_hd__buf_1 _2543_ (
    .A(_0177_),
    .X(_0242_)
  );
  sky130_fd_sc_hd__or3_2 _2544_ (
    .A(_0123_),
    .B(_0242_),
    .C(_0166_),
    .X(_0243_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2545_ (
    .A1(_0113_),
    .A2(_0237_),
    .B1(_0238_),
    .C1(_0241_),
    .D1(_0243_),
    .Y(_0244_)
  );
  sky130_fd_sc_hd__or4_2 _2546_ (
    .A(_0214_),
    .B(_0223_),
    .C(_0234_),
    .D(_0244_),
    .X(_0245_)
  );
  sky130_fd_sc_hd__or4_2 _2547_ (
    .A(_0161_),
    .B(_0181_),
    .C(_0203_),
    .D(_0245_),
    .X(_0246_)
  );
  sky130_fd_sc_hd__buf_1 _2548_ (
    .A(_0246_),
    .X(\g_bit[31].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _2549_ (
    .A1(\g_bit[0].g_word[30].r_bit.Q ),
    .A2(_0023_),
    .A3(_0025_),
    .B1(_0030_),
    .B2(\g_bit[0].g_word[28].r_bit.Q ),
    .X(_0247_)
  );
  sky130_fd_sc_hd__a221o_2 _2550_ (
    .A1(\g_bit[0].g_word[4].r_bit.Q ),
    .A2(_0014_),
    .B1(_0021_),
    .B2(\g_bit[0].g_word[26].r_bit.Q ),
    .C1(_0247_),
    .X(_0248_)
  );
  sky130_fd_sc_hd__a22o_2 _2551_ (
    .A1(\g_bit[0].g_word[5].r_bit.Q ),
    .A2(_0043_),
    .B1(_0050_),
    .B2(\g_bit[0].g_word[2].r_bit.Q ),
    .X(_0249_)
  );
  sky130_fd_sc_hd__a221o_2 _2552_ (
    .A1(\g_bit[0].g_word[25].r_bit.Q ),
    .A2(_0035_),
    .B1(_0039_),
    .B2(\g_bit[0].g_word[31].r_bit.Q ),
    .C1(_0249_),
    .X(_0250_)
  );
  sky130_fd_sc_hd__a22o_2 _2553_ (
    .A1(\g_bit[0].g_word[13].r_bit.Q ),
    .A2(_0054_),
    .B1(_0057_),
    .B2(\g_bit[0].g_word[15].r_bit.Q ),
    .X(_0251_)
  );
  sky130_fd_sc_hd__a22o_2 _2554_ (
    .A1(\g_bit[0].g_word[11].r_bit.Q ),
    .A2(_0060_),
    .B1(_0062_),
    .B2(\g_bit[0].g_word[20].r_bit.Q ),
    .X(_0252_)
  );
  sky130_fd_sc_hd__a22o_2 _2555_ (
    .A1(\g_bit[0].g_word[19].r_bit.Q ),
    .A2(_0065_),
    .B1(_0067_),
    .B2(\g_bit[0].g_word[21].r_bit.Q ),
    .X(_0253_)
  );
  sky130_fd_sc_hd__a22o_2 _2556_ (
    .A1(\g_bit[0].g_word[17].r_bit.Q ),
    .A2(_0070_),
    .B1(_0072_),
    .B2(\g_bit[0].g_word[12].r_bit.Q ),
    .X(_0254_)
  );
  sky130_fd_sc_hd__or4_2 _2557_ (
    .A(_0251_),
    .B(_0252_),
    .C(_0253_),
    .D(_0254_),
    .X(_0255_)
  );
  sky130_fd_sc_hd__inv_2 _2558_ (
    .A(\g_bit[0].g_word[7].r_bit.Q ),
    .Y(_0256_)
  );
  sky130_fd_sc_hd__nor3_2 _2559_ (
    .A(_0256_),
    .B(_0082_),
    .C(_0004_),
    .Y(_0257_)
  );
  sky130_fd_sc_hd__inv_2 _2560_ (
    .A(\g_bit[0].g_word[3].r_bit.Q ),
    .Y(_0258_)
  );
  sky130_fd_sc_hd__nor3_2 _2561_ (
    .A(_0258_),
    .B(_0085_),
    .C(_0086_),
    .Y(_0259_)
  );
  sky130_fd_sc_hd__buf_1 _2562_ (
    .A(_0077_),
    .X(_0260_)
  );
  sky130_fd_sc_hd__buf_1 _2563_ (
    .A(_0078_),
    .X(_0261_)
  );
  sky130_fd_sc_hd__and3_2 _2564_ (
    .A(\g_bit[0].g_word[24].r_bit.Q ),
    .B(_0260_),
    .C(_0261_),
    .X(_0262_)
  );
  sky130_fd_sc_hd__a2111o_2 _2565_ (
    .A1(\g_bit[0].g_word[29].r_bit.Q ),
    .A2(_0076_),
    .B1(_0257_),
    .C1(_0259_),
    .D1(_0262_),
    .X(_0263_)
  );
  sky130_fd_sc_hd__and3_2 _2566_ (
    .A(\g_bit[0].g_word[27].r_bit.Q ),
    .B(_0094_),
    .C(_0095_),
    .X(_0264_)
  );
  sky130_fd_sc_hd__a221o_2 _2567_ (
    .A1(\g_bit[0].g_word[6].r_bit.Q ),
    .A2(_0090_),
    .B1(_0092_),
    .B2(\g_bit[0].g_word[1].r_bit.Q ),
    .C1(_0264_),
    .X(_0265_)
  );
  sky130_fd_sc_hd__inv_2 _2568_ (
    .A(\g_bit[0].g_word[23].r_bit.Q ),
    .Y(_0266_)
  );
  sky130_fd_sc_hd__inv_2 _2569_ (
    .A(\g_bit[0].g_word[10].r_bit.Q ),
    .Y(_0267_)
  );
  sky130_fd_sc_hd__or3_2 _2570_ (
    .A(_0267_),
    .B(_0103_),
    .C(_0107_),
    .X(_0268_)
  );
  sky130_fd_sc_hd__inv_2 _2571_ (
    .A(\g_bit[0].g_word[9].r_bit.Q ),
    .Y(_0269_)
  );
  sky130_fd_sc_hd__or3_2 _2572_ (
    .A(_0269_),
    .B(_0106_),
    .C(_0110_),
    .X(_0270_)
  );
  sky130_fd_sc_hd__inv_2 _2573_ (
    .A(\g_bit[0].g_word[8].r_bit.Q ),
    .Y(_0271_)
  );
  sky130_fd_sc_hd__or3_2 _2574_ (
    .A(_0271_),
    .B(_0017_),
    .C(_0012_),
    .X(_0272_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2575_ (
    .A1(_0266_),
    .A2(_0101_),
    .B1(_0268_),
    .C1(_0270_),
    .D1(_0272_),
    .Y(_0273_)
  );
  sky130_fd_sc_hd__inv_2 _2576_ (
    .A(\g_bit[0].g_word[22].r_bit.Q ),
    .Y(_0274_)
  );
  sky130_fd_sc_hd__inv_2 _2577_ (
    .A(\g_bit[0].g_word[16].r_bit.Q ),
    .Y(_0275_)
  );
  sky130_fd_sc_hd__or3_2 _2578_ (
    .A(_0275_),
    .B(_0118_),
    .C(_0121_),
    .X(_0276_)
  );
  sky130_fd_sc_hd__inv_2 _2579_ (
    .A(\g_bit[0].g_word[14].r_bit.Q ),
    .Y(_0277_)
  );
  sky130_fd_sc_hd__or3_2 _2580_ (
    .A(_0277_),
    .B(_0124_),
    .C(_0037_),
    .X(_0278_)
  );
  sky130_fd_sc_hd__inv_2 _2581_ (
    .A(\g_bit[0].g_word[18].r_bit.Q ),
    .Y(_0279_)
  );
  sky130_fd_sc_hd__buf_1 _2582_ (
    .A(_0046_),
    .X(_0280_)
  );
  sky130_fd_sc_hd__or3_2 _2583_ (
    .A(_0279_),
    .B(_0280_),
    .C(_0019_),
    .X(_0281_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2584_ (
    .A1(_0274_),
    .A2(_0116_),
    .B1(_0276_),
    .C1(_0278_),
    .D1(_0281_),
    .Y(_0282_)
  );
  sky130_fd_sc_hd__or4_2 _2585_ (
    .A(_0263_),
    .B(_0265_),
    .C(_0273_),
    .D(_0282_),
    .X(_0283_)
  );
  sky130_fd_sc_hd__or4_2 _2586_ (
    .A(_0248_),
    .B(_0250_),
    .C(_0255_),
    .D(_0283_),
    .X(_0284_)
  );
  sky130_fd_sc_hd__buf_1 _2587_ (
    .A(_0284_),
    .X(\g_bit[0].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _2588_ (
    .A1(\g_bit[0].g_word[30].r_bit.Q ),
    .A2(_0152_),
    .A3(_0154_),
    .B1(_0159_),
    .B2(\g_bit[0].g_word[28].r_bit.Q ),
    .X(_0285_)
  );
  sky130_fd_sc_hd__a221o_2 _2589_ (
    .A1(\g_bit[0].g_word[4].r_bit.Q ),
    .A2(_0143_),
    .B1(_0150_),
    .B2(\g_bit[0].g_word[26].r_bit.Q ),
    .C1(_0285_),
    .X(_0286_)
  );
  sky130_fd_sc_hd__a22o_2 _2590_ (
    .A1(\g_bit[0].g_word[5].r_bit.Q ),
    .A2(_0172_),
    .B1(_0179_),
    .B2(\g_bit[0].g_word[2].r_bit.Q ),
    .X(_0287_)
  );
  sky130_fd_sc_hd__a221o_2 _2591_ (
    .A1(\g_bit[0].g_word[25].r_bit.Q ),
    .A2(_0164_),
    .B1(_0168_),
    .B2(\g_bit[0].g_word[31].r_bit.Q ),
    .C1(_0287_),
    .X(_0288_)
  );
  sky130_fd_sc_hd__a22o_2 _2592_ (
    .A1(\g_bit[0].g_word[13].r_bit.Q ),
    .A2(_0183_),
    .B1(_0186_),
    .B2(\g_bit[0].g_word[15].r_bit.Q ),
    .X(_0289_)
  );
  sky130_fd_sc_hd__a22o_2 _2593_ (
    .A1(\g_bit[0].g_word[20].r_bit.Q ),
    .A2(_0189_),
    .B1(_0191_),
    .B2(\g_bit[0].g_word[11].r_bit.Q ),
    .X(_0290_)
  );
  sky130_fd_sc_hd__a22o_2 _2594_ (
    .A1(\g_bit[0].g_word[19].r_bit.Q ),
    .A2(_0194_),
    .B1(_0196_),
    .B2(\g_bit[0].g_word[21].r_bit.Q ),
    .X(_0291_)
  );
  sky130_fd_sc_hd__a22o_2 _2595_ (
    .A1(\g_bit[0].g_word[17].r_bit.Q ),
    .A2(_0199_),
    .B1(_0201_),
    .B2(\g_bit[0].g_word[12].r_bit.Q ),
    .X(_0292_)
  );
  sky130_fd_sc_hd__or4_2 _2596_ (
    .A(_0289_),
    .B(_0290_),
    .C(_0291_),
    .D(_0292_),
    .X(_0293_)
  );
  sky130_fd_sc_hd__buf_1 _2597_ (
    .A(_0209_),
    .X(_0294_)
  );
  sky130_fd_sc_hd__nor3_2 _2598_ (
    .A(_0256_),
    .B(_0133_),
    .C(_0294_),
    .Y(_0295_)
  );
  sky130_fd_sc_hd__nor3_2 _2599_ (
    .A(_0258_),
    .B(_0212_),
    .C(_0210_),
    .Y(_0296_)
  );
  sky130_fd_sc_hd__buf_1 _2600_ (
    .A(_0206_),
    .X(_0297_)
  );
  sky130_fd_sc_hd__buf_1 _2601_ (
    .A(_0207_),
    .X(_0298_)
  );
  sky130_fd_sc_hd__and3_2 _2602_ (
    .A(\g_bit[0].g_word[24].r_bit.Q ),
    .B(_0297_),
    .C(_0298_),
    .X(_0299_)
  );
  sky130_fd_sc_hd__a2111o_2 _2603_ (
    .A1(\g_bit[0].g_word[29].r_bit.Q ),
    .A2(_0205_),
    .B1(_0295_),
    .C1(_0296_),
    .D1(_0299_),
    .X(_0300_)
  );
  sky130_fd_sc_hd__and3_2 _2604_ (
    .A(\g_bit[0].g_word[27].r_bit.Q ),
    .B(_0220_),
    .C(_0221_),
    .X(_0301_)
  );
  sky130_fd_sc_hd__a221o_2 _2605_ (
    .A1(\g_bit[0].g_word[6].r_bit.Q ),
    .A2(_0216_),
    .B1(_0218_),
    .B2(\g_bit[0].g_word[1].r_bit.Q ),
    .C1(_0301_),
    .X(_0302_)
  );
  sky130_fd_sc_hd__or3_2 _2606_ (
    .A(_0267_),
    .B(_0227_),
    .C(_0230_),
    .X(_0303_)
  );
  sky130_fd_sc_hd__or3_2 _2607_ (
    .A(_0269_),
    .B(_0229_),
    .C(_0232_),
    .X(_0304_)
  );
  sky130_fd_sc_hd__or3_2 _2608_ (
    .A(_0271_),
    .B(_0146_),
    .C(_0141_),
    .X(_0305_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2609_ (
    .A1(_0266_),
    .A2(_0226_),
    .B1(_0303_),
    .C1(_0304_),
    .D1(_0305_),
    .Y(_0306_)
  );
  sky130_fd_sc_hd__or3_2 _2610_ (
    .A(_0275_),
    .B(_0239_),
    .C(_0240_),
    .X(_0307_)
  );
  sky130_fd_sc_hd__or3_2 _2611_ (
    .A(_0277_),
    .B(_0242_),
    .C(_0166_),
    .X(_0308_)
  );
  sky130_fd_sc_hd__buf_1 _2612_ (
    .A(_0175_),
    .X(_0309_)
  );
  sky130_fd_sc_hd__or3_2 _2613_ (
    .A(_0279_),
    .B(_0309_),
    .C(_0148_),
    .X(_0310_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2614_ (
    .A1(_0274_),
    .A2(_0237_),
    .B1(_0307_),
    .C1(_0308_),
    .D1(_0310_),
    .Y(_0311_)
  );
  sky130_fd_sc_hd__or4_2 _2615_ (
    .A(_0300_),
    .B(_0302_),
    .C(_0306_),
    .D(_0311_),
    .X(_0312_)
  );
  sky130_fd_sc_hd__or4_2 _2616_ (
    .A(_0286_),
    .B(_0288_),
    .C(_0293_),
    .D(_0312_),
    .X(_0313_)
  );
  sky130_fd_sc_hd__buf_1 _2617_ (
    .A(_0313_),
    .X(\g_bit[0].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _2618_ (
    .A1(\g_bit[1].g_word[30].r_bit.Q ),
    .A2(_0023_),
    .A3(_0025_),
    .B1(_0030_),
    .B2(\g_bit[1].g_word[28].r_bit.Q ),
    .X(_0314_)
  );
  sky130_fd_sc_hd__a221o_2 _2619_ (
    .A1(\g_bit[1].g_word[4].r_bit.Q ),
    .A2(_0014_),
    .B1(_0021_),
    .B2(\g_bit[1].g_word[26].r_bit.Q ),
    .C1(_0314_),
    .X(_0315_)
  );
  sky130_fd_sc_hd__a22o_2 _2620_ (
    .A1(\g_bit[1].g_word[5].r_bit.Q ),
    .A2(_0043_),
    .B1(_0050_),
    .B2(\g_bit[1].g_word[2].r_bit.Q ),
    .X(_0316_)
  );
  sky130_fd_sc_hd__a221o_2 _2621_ (
    .A1(\g_bit[1].g_word[25].r_bit.Q ),
    .A2(_0035_),
    .B1(_0039_),
    .B2(\g_bit[1].g_word[31].r_bit.Q ),
    .C1(_0316_),
    .X(_0317_)
  );
  sky130_fd_sc_hd__a22o_2 _2622_ (
    .A1(\g_bit[1].g_word[13].r_bit.Q ),
    .A2(_0054_),
    .B1(_0057_),
    .B2(\g_bit[1].g_word[15].r_bit.Q ),
    .X(_0318_)
  );
  sky130_fd_sc_hd__a22o_2 _2623_ (
    .A1(\g_bit[1].g_word[11].r_bit.Q ),
    .A2(_0060_),
    .B1(_0062_),
    .B2(\g_bit[1].g_word[20].r_bit.Q ),
    .X(_0319_)
  );
  sky130_fd_sc_hd__a22o_2 _2624_ (
    .A1(\g_bit[1].g_word[19].r_bit.Q ),
    .A2(_0065_),
    .B1(_0067_),
    .B2(\g_bit[1].g_word[21].r_bit.Q ),
    .X(_0320_)
  );
  sky130_fd_sc_hd__a22o_2 _2625_ (
    .A1(\g_bit[1].g_word[17].r_bit.Q ),
    .A2(_0070_),
    .B1(_0072_),
    .B2(\g_bit[1].g_word[12].r_bit.Q ),
    .X(_0321_)
  );
  sky130_fd_sc_hd__or4_2 _2626_ (
    .A(_0318_),
    .B(_0319_),
    .C(_0320_),
    .D(_0321_),
    .X(_0322_)
  );
  sky130_fd_sc_hd__inv_2 _2627_ (
    .A(\g_bit[1].g_word[7].r_bit.Q ),
    .Y(_0323_)
  );
  sky130_fd_sc_hd__nor3_2 _2628_ (
    .A(_0323_),
    .B(_0082_),
    .C(_0004_),
    .Y(_0324_)
  );
  sky130_fd_sc_hd__inv_2 _2629_ (
    .A(\g_bit[1].g_word[3].r_bit.Q ),
    .Y(_0325_)
  );
  sky130_fd_sc_hd__nor3_2 _2630_ (
    .A(_0325_),
    .B(_0085_),
    .C(_0086_),
    .Y(_0326_)
  );
  sky130_fd_sc_hd__and3_2 _2631_ (
    .A(\g_bit[1].g_word[24].r_bit.Q ),
    .B(_0260_),
    .C(_0261_),
    .X(_0327_)
  );
  sky130_fd_sc_hd__a2111o_2 _2632_ (
    .A1(\g_bit[1].g_word[29].r_bit.Q ),
    .A2(_0076_),
    .B1(_0324_),
    .C1(_0326_),
    .D1(_0327_),
    .X(_0328_)
  );
  sky130_fd_sc_hd__and3_2 _2633_ (
    .A(\g_bit[1].g_word[27].r_bit.Q ),
    .B(_0094_),
    .C(_0095_),
    .X(_0329_)
  );
  sky130_fd_sc_hd__a221o_2 _2634_ (
    .A1(\g_bit[1].g_word[6].r_bit.Q ),
    .A2(_0090_),
    .B1(_0092_),
    .B2(\g_bit[1].g_word[1].r_bit.Q ),
    .C1(_0329_),
    .X(_0330_)
  );
  sky130_fd_sc_hd__inv_2 _2635_ (
    .A(\g_bit[1].g_word[23].r_bit.Q ),
    .Y(_0331_)
  );
  sky130_fd_sc_hd__inv_2 _2636_ (
    .A(\g_bit[1].g_word[10].r_bit.Q ),
    .Y(_0332_)
  );
  sky130_fd_sc_hd__or3_2 _2637_ (
    .A(_0332_),
    .B(_0103_),
    .C(_0107_),
    .X(_0333_)
  );
  sky130_fd_sc_hd__inv_2 _2638_ (
    .A(\g_bit[1].g_word[9].r_bit.Q ),
    .Y(_0334_)
  );
  sky130_fd_sc_hd__or3_2 _2639_ (
    .A(_0334_),
    .B(_0106_),
    .C(_0110_),
    .X(_0335_)
  );
  sky130_fd_sc_hd__inv_2 _2640_ (
    .A(\g_bit[1].g_word[8].r_bit.Q ),
    .Y(_0336_)
  );
  sky130_fd_sc_hd__or3_2 _2641_ (
    .A(_0336_),
    .B(_0017_),
    .C(_0012_),
    .X(_0337_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2642_ (
    .A1(_0331_),
    .A2(_0101_),
    .B1(_0333_),
    .C1(_0335_),
    .D1(_0337_),
    .Y(_0338_)
  );
  sky130_fd_sc_hd__inv_2 _2643_ (
    .A(\g_bit[1].g_word[22].r_bit.Q ),
    .Y(_0339_)
  );
  sky130_fd_sc_hd__inv_2 _2644_ (
    .A(\g_bit[1].g_word[16].r_bit.Q ),
    .Y(_0340_)
  );
  sky130_fd_sc_hd__or3_2 _2645_ (
    .A(_0340_),
    .B(_0118_),
    .C(_0121_),
    .X(_0341_)
  );
  sky130_fd_sc_hd__inv_2 _2646_ (
    .A(\g_bit[1].g_word[14].r_bit.Q ),
    .Y(_0342_)
  );
  sky130_fd_sc_hd__or3_2 _2647_ (
    .A(_0342_),
    .B(_0124_),
    .C(_0037_),
    .X(_0343_)
  );
  sky130_fd_sc_hd__inv_2 _2648_ (
    .A(\g_bit[1].g_word[18].r_bit.Q ),
    .Y(_0344_)
  );
  sky130_fd_sc_hd__or3_2 _2649_ (
    .A(_0344_),
    .B(_0280_),
    .C(_0019_),
    .X(_0345_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2650_ (
    .A1(_0339_),
    .A2(_0116_),
    .B1(_0341_),
    .C1(_0343_),
    .D1(_0345_),
    .Y(_0346_)
  );
  sky130_fd_sc_hd__or4_2 _2651_ (
    .A(_0328_),
    .B(_0330_),
    .C(_0338_),
    .D(_0346_),
    .X(_0347_)
  );
  sky130_fd_sc_hd__or4_2 _2652_ (
    .A(_0315_),
    .B(_0317_),
    .C(_0322_),
    .D(_0347_),
    .X(_0348_)
  );
  sky130_fd_sc_hd__buf_1 _2653_ (
    .A(_0348_),
    .X(\g_bit[1].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _2654_ (
    .A1(\g_bit[1].g_word[30].r_bit.Q ),
    .A2(_0152_),
    .A3(_0154_),
    .B1(_0159_),
    .B2(\g_bit[1].g_word[28].r_bit.Q ),
    .X(_0349_)
  );
  sky130_fd_sc_hd__a221o_2 _2655_ (
    .A1(\g_bit[1].g_word[4].r_bit.Q ),
    .A2(_0143_),
    .B1(_0150_),
    .B2(\g_bit[1].g_word[26].r_bit.Q ),
    .C1(_0349_),
    .X(_0350_)
  );
  sky130_fd_sc_hd__a22o_2 _2656_ (
    .A1(\g_bit[1].g_word[5].r_bit.Q ),
    .A2(_0172_),
    .B1(_0179_),
    .B2(\g_bit[1].g_word[2].r_bit.Q ),
    .X(_0351_)
  );
  sky130_fd_sc_hd__a221o_2 _2657_ (
    .A1(\g_bit[1].g_word[25].r_bit.Q ),
    .A2(_0164_),
    .B1(_0168_),
    .B2(\g_bit[1].g_word[31].r_bit.Q ),
    .C1(_0351_),
    .X(_0352_)
  );
  sky130_fd_sc_hd__a22o_2 _2658_ (
    .A1(\g_bit[1].g_word[13].r_bit.Q ),
    .A2(_0183_),
    .B1(_0186_),
    .B2(\g_bit[1].g_word[15].r_bit.Q ),
    .X(_0353_)
  );
  sky130_fd_sc_hd__a22o_2 _2659_ (
    .A1(\g_bit[1].g_word[20].r_bit.Q ),
    .A2(_0189_),
    .B1(_0191_),
    .B2(\g_bit[1].g_word[11].r_bit.Q ),
    .X(_0354_)
  );
  sky130_fd_sc_hd__a22o_2 _2660_ (
    .A1(\g_bit[1].g_word[19].r_bit.Q ),
    .A2(_0194_),
    .B1(_0196_),
    .B2(\g_bit[1].g_word[21].r_bit.Q ),
    .X(_0355_)
  );
  sky130_fd_sc_hd__a22o_2 _2661_ (
    .A1(\g_bit[1].g_word[17].r_bit.Q ),
    .A2(_0199_),
    .B1(_0201_),
    .B2(\g_bit[1].g_word[12].r_bit.Q ),
    .X(_0356_)
  );
  sky130_fd_sc_hd__or4_2 _2662_ (
    .A(_0353_),
    .B(_0354_),
    .C(_0355_),
    .D(_0356_),
    .X(_0357_)
  );
  sky130_fd_sc_hd__nor3_2 _2663_ (
    .A(_0323_),
    .B(_0133_),
    .C(_0294_),
    .Y(_0358_)
  );
  sky130_fd_sc_hd__nor3_2 _2664_ (
    .A(_0325_),
    .B(_0212_),
    .C(_0210_),
    .Y(_0359_)
  );
  sky130_fd_sc_hd__and3_2 _2665_ (
    .A(\g_bit[1].g_word[24].r_bit.Q ),
    .B(_0297_),
    .C(_0298_),
    .X(_0360_)
  );
  sky130_fd_sc_hd__a2111o_2 _2666_ (
    .A1(\g_bit[1].g_word[29].r_bit.Q ),
    .A2(_0205_),
    .B1(_0358_),
    .C1(_0359_),
    .D1(_0360_),
    .X(_0361_)
  );
  sky130_fd_sc_hd__and3_2 _2667_ (
    .A(\g_bit[1].g_word[27].r_bit.Q ),
    .B(_0220_),
    .C(_0221_),
    .X(_0362_)
  );
  sky130_fd_sc_hd__a221o_2 _2668_ (
    .A1(\g_bit[1].g_word[6].r_bit.Q ),
    .A2(_0216_),
    .B1(_0218_),
    .B2(\g_bit[1].g_word[1].r_bit.Q ),
    .C1(_0362_),
    .X(_0363_)
  );
  sky130_fd_sc_hd__or3_2 _2669_ (
    .A(_0332_),
    .B(_0227_),
    .C(_0230_),
    .X(_0364_)
  );
  sky130_fd_sc_hd__or3_2 _2670_ (
    .A(_0334_),
    .B(_0229_),
    .C(_0232_),
    .X(_0365_)
  );
  sky130_fd_sc_hd__or3_2 _2671_ (
    .A(_0336_),
    .B(_0146_),
    .C(_0141_),
    .X(_0366_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2672_ (
    .A1(_0331_),
    .A2(_0226_),
    .B1(_0364_),
    .C1(_0365_),
    .D1(_0366_),
    .Y(_0367_)
  );
  sky130_fd_sc_hd__or3_2 _2673_ (
    .A(_0340_),
    .B(_0239_),
    .C(_0240_),
    .X(_0368_)
  );
  sky130_fd_sc_hd__or3_2 _2674_ (
    .A(_0342_),
    .B(_0242_),
    .C(_0166_),
    .X(_0369_)
  );
  sky130_fd_sc_hd__or3_2 _2675_ (
    .A(_0344_),
    .B(_0309_),
    .C(_0148_),
    .X(_0370_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2676_ (
    .A1(_0339_),
    .A2(_0237_),
    .B1(_0368_),
    .C1(_0369_),
    .D1(_0370_),
    .Y(_0371_)
  );
  sky130_fd_sc_hd__or4_2 _2677_ (
    .A(_0361_),
    .B(_0363_),
    .C(_0367_),
    .D(_0371_),
    .X(_0372_)
  );
  sky130_fd_sc_hd__or4_2 _2678_ (
    .A(_0350_),
    .B(_0352_),
    .C(_0357_),
    .D(_0372_),
    .X(_0373_)
  );
  sky130_fd_sc_hd__buf_1 _2679_ (
    .A(_0373_),
    .X(\g_bit[1].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _2680_ (
    .A1(\g_bit[2].g_word[30].r_bit.Q ),
    .A2(_0023_),
    .A3(_0025_),
    .B1(_0030_),
    .B2(\g_bit[2].g_word[28].r_bit.Q ),
    .X(_0374_)
  );
  sky130_fd_sc_hd__a221o_2 _2681_ (
    .A1(\g_bit[2].g_word[4].r_bit.Q ),
    .A2(_0014_),
    .B1(_0021_),
    .B2(\g_bit[2].g_word[26].r_bit.Q ),
    .C1(_0374_),
    .X(_0375_)
  );
  sky130_fd_sc_hd__a22o_2 _2682_ (
    .A1(\g_bit[2].g_word[5].r_bit.Q ),
    .A2(_0043_),
    .B1(_0050_),
    .B2(\g_bit[2].g_word[2].r_bit.Q ),
    .X(_0376_)
  );
  sky130_fd_sc_hd__a221o_2 _2683_ (
    .A1(\g_bit[2].g_word[25].r_bit.Q ),
    .A2(_0035_),
    .B1(_0039_),
    .B2(\g_bit[2].g_word[31].r_bit.Q ),
    .C1(_0376_),
    .X(_0377_)
  );
  sky130_fd_sc_hd__a22o_2 _2684_ (
    .A1(\g_bit[2].g_word[13].r_bit.Q ),
    .A2(_0054_),
    .B1(_0057_),
    .B2(\g_bit[2].g_word[15].r_bit.Q ),
    .X(_0378_)
  );
  sky130_fd_sc_hd__a22o_2 _2685_ (
    .A1(\g_bit[2].g_word[11].r_bit.Q ),
    .A2(_0060_),
    .B1(_0062_),
    .B2(\g_bit[2].g_word[20].r_bit.Q ),
    .X(_0379_)
  );
  sky130_fd_sc_hd__a22o_2 _2686_ (
    .A1(\g_bit[2].g_word[19].r_bit.Q ),
    .A2(_0065_),
    .B1(_0067_),
    .B2(\g_bit[2].g_word[21].r_bit.Q ),
    .X(_0380_)
  );
  sky130_fd_sc_hd__a22o_2 _2687_ (
    .A1(\g_bit[2].g_word[17].r_bit.Q ),
    .A2(_0070_),
    .B1(_0072_),
    .B2(\g_bit[2].g_word[12].r_bit.Q ),
    .X(_0381_)
  );
  sky130_fd_sc_hd__or4_2 _2688_ (
    .A(_0378_),
    .B(_0379_),
    .C(_0380_),
    .D(_0381_),
    .X(_0382_)
  );
  sky130_fd_sc_hd__inv_2 _2689_ (
    .A(\g_bit[2].g_word[7].r_bit.Q ),
    .Y(_0383_)
  );
  sky130_fd_sc_hd__nor3_2 _2690_ (
    .A(_0383_),
    .B(_0082_),
    .C(_0004_),
    .Y(_0384_)
  );
  sky130_fd_sc_hd__inv_2 _2691_ (
    .A(\g_bit[2].g_word[3].r_bit.Q ),
    .Y(_0385_)
  );
  sky130_fd_sc_hd__nor3_2 _2692_ (
    .A(_0385_),
    .B(_0085_),
    .C(_0086_),
    .Y(_0386_)
  );
  sky130_fd_sc_hd__and3_2 _2693_ (
    .A(\g_bit[2].g_word[24].r_bit.Q ),
    .B(_0260_),
    .C(_0261_),
    .X(_0387_)
  );
  sky130_fd_sc_hd__a2111o_2 _2694_ (
    .A1(\g_bit[2].g_word[29].r_bit.Q ),
    .A2(_0076_),
    .B1(_0384_),
    .C1(_0386_),
    .D1(_0387_),
    .X(_0388_)
  );
  sky130_fd_sc_hd__and3_2 _2695_ (
    .A(\g_bit[2].g_word[27].r_bit.Q ),
    .B(_0094_),
    .C(_0095_),
    .X(_0389_)
  );
  sky130_fd_sc_hd__a221o_2 _2696_ (
    .A1(\g_bit[2].g_word[6].r_bit.Q ),
    .A2(_0090_),
    .B1(_0092_),
    .B2(\g_bit[2].g_word[1].r_bit.Q ),
    .C1(_0389_),
    .X(_0390_)
  );
  sky130_fd_sc_hd__inv_2 _2697_ (
    .A(\g_bit[2].g_word[23].r_bit.Q ),
    .Y(_0391_)
  );
  sky130_fd_sc_hd__inv_2 _2698_ (
    .A(\g_bit[2].g_word[10].r_bit.Q ),
    .Y(_0392_)
  );
  sky130_fd_sc_hd__or3_2 _2699_ (
    .A(_0392_),
    .B(_0103_),
    .C(_0107_),
    .X(_0393_)
  );
  sky130_fd_sc_hd__inv_2 _2700_ (
    .A(\g_bit[2].g_word[9].r_bit.Q ),
    .Y(_0394_)
  );
  sky130_fd_sc_hd__or3_2 _2701_ (
    .A(_0394_),
    .B(_0106_),
    .C(_0110_),
    .X(_0395_)
  );
  sky130_fd_sc_hd__inv_2 _2702_ (
    .A(\g_bit[2].g_word[8].r_bit.Q ),
    .Y(_0396_)
  );
  sky130_fd_sc_hd__or3_2 _2703_ (
    .A(_0396_),
    .B(_0017_),
    .C(_0012_),
    .X(_0397_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2704_ (
    .A1(_0391_),
    .A2(_0101_),
    .B1(_0393_),
    .C1(_0395_),
    .D1(_0397_),
    .Y(_0398_)
  );
  sky130_fd_sc_hd__inv_2 _2705_ (
    .A(\g_bit[2].g_word[22].r_bit.Q ),
    .Y(_0399_)
  );
  sky130_fd_sc_hd__inv_2 _2706_ (
    .A(\g_bit[2].g_word[16].r_bit.Q ),
    .Y(_0400_)
  );
  sky130_fd_sc_hd__or3_2 _2707_ (
    .A(_0400_),
    .B(_0118_),
    .C(_0121_),
    .X(_0401_)
  );
  sky130_fd_sc_hd__inv_2 _2708_ (
    .A(\g_bit[2].g_word[14].r_bit.Q ),
    .Y(_0402_)
  );
  sky130_fd_sc_hd__or3_2 _2709_ (
    .A(_0402_),
    .B(_0124_),
    .C(_0037_),
    .X(_0403_)
  );
  sky130_fd_sc_hd__inv_2 _2710_ (
    .A(\g_bit[2].g_word[18].r_bit.Q ),
    .Y(_0404_)
  );
  sky130_fd_sc_hd__or3_2 _2711_ (
    .A(_0404_),
    .B(_0280_),
    .C(_0019_),
    .X(_0405_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2712_ (
    .A1(_0399_),
    .A2(_0116_),
    .B1(_0401_),
    .C1(_0403_),
    .D1(_0405_),
    .Y(_0406_)
  );
  sky130_fd_sc_hd__or4_2 _2713_ (
    .A(_0388_),
    .B(_0390_),
    .C(_0398_),
    .D(_0406_),
    .X(_0407_)
  );
  sky130_fd_sc_hd__or4_2 _2714_ (
    .A(_0375_),
    .B(_0377_),
    .C(_0382_),
    .D(_0407_),
    .X(_0408_)
  );
  sky130_fd_sc_hd__buf_1 _2715_ (
    .A(_0408_),
    .X(\g_bit[2].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _2716_ (
    .A1(\g_bit[2].g_word[30].r_bit.Q ),
    .A2(_0152_),
    .A3(_0154_),
    .B1(_0159_),
    .B2(\g_bit[2].g_word[28].r_bit.Q ),
    .X(_0409_)
  );
  sky130_fd_sc_hd__a221o_2 _2717_ (
    .A1(\g_bit[2].g_word[4].r_bit.Q ),
    .A2(_0143_),
    .B1(_0150_),
    .B2(\g_bit[2].g_word[26].r_bit.Q ),
    .C1(_0409_),
    .X(_0410_)
  );
  sky130_fd_sc_hd__a22o_2 _2718_ (
    .A1(\g_bit[2].g_word[5].r_bit.Q ),
    .A2(_0172_),
    .B1(_0179_),
    .B2(\g_bit[2].g_word[2].r_bit.Q ),
    .X(_0411_)
  );
  sky130_fd_sc_hd__a221o_2 _2719_ (
    .A1(\g_bit[2].g_word[25].r_bit.Q ),
    .A2(_0164_),
    .B1(_0168_),
    .B2(\g_bit[2].g_word[31].r_bit.Q ),
    .C1(_0411_),
    .X(_0412_)
  );
  sky130_fd_sc_hd__a22o_2 _2720_ (
    .A1(\g_bit[2].g_word[13].r_bit.Q ),
    .A2(_0183_),
    .B1(_0186_),
    .B2(\g_bit[2].g_word[15].r_bit.Q ),
    .X(_0413_)
  );
  sky130_fd_sc_hd__a22o_2 _2721_ (
    .A1(\g_bit[2].g_word[20].r_bit.Q ),
    .A2(_0189_),
    .B1(_0191_),
    .B2(\g_bit[2].g_word[11].r_bit.Q ),
    .X(_0414_)
  );
  sky130_fd_sc_hd__a22o_2 _2722_ (
    .A1(\g_bit[2].g_word[19].r_bit.Q ),
    .A2(_0194_),
    .B1(_0196_),
    .B2(\g_bit[2].g_word[21].r_bit.Q ),
    .X(_0415_)
  );
  sky130_fd_sc_hd__a22o_2 _2723_ (
    .A1(\g_bit[2].g_word[17].r_bit.Q ),
    .A2(_0199_),
    .B1(_0201_),
    .B2(\g_bit[2].g_word[12].r_bit.Q ),
    .X(_0416_)
  );
  sky130_fd_sc_hd__or4_2 _2724_ (
    .A(_0413_),
    .B(_0414_),
    .C(_0415_),
    .D(_0416_),
    .X(_0417_)
  );
  sky130_fd_sc_hd__nor3_2 _2725_ (
    .A(_0383_),
    .B(_0133_),
    .C(_0294_),
    .Y(_0418_)
  );
  sky130_fd_sc_hd__nor3_2 _2726_ (
    .A(_0385_),
    .B(_0212_),
    .C(_0210_),
    .Y(_0419_)
  );
  sky130_fd_sc_hd__and3_2 _2727_ (
    .A(\g_bit[2].g_word[24].r_bit.Q ),
    .B(_0297_),
    .C(_0298_),
    .X(_0420_)
  );
  sky130_fd_sc_hd__a2111o_2 _2728_ (
    .A1(\g_bit[2].g_word[29].r_bit.Q ),
    .A2(_0205_),
    .B1(_0418_),
    .C1(_0419_),
    .D1(_0420_),
    .X(_0421_)
  );
  sky130_fd_sc_hd__and3_2 _2729_ (
    .A(\g_bit[2].g_word[27].r_bit.Q ),
    .B(_0220_),
    .C(_0221_),
    .X(_0422_)
  );
  sky130_fd_sc_hd__a221o_2 _2730_ (
    .A1(\g_bit[2].g_word[6].r_bit.Q ),
    .A2(_0216_),
    .B1(_0218_),
    .B2(\g_bit[2].g_word[1].r_bit.Q ),
    .C1(_0422_),
    .X(_0423_)
  );
  sky130_fd_sc_hd__or3_2 _2731_ (
    .A(_0392_),
    .B(_0227_),
    .C(_0230_),
    .X(_0424_)
  );
  sky130_fd_sc_hd__or3_2 _2732_ (
    .A(_0394_),
    .B(_0229_),
    .C(_0232_),
    .X(_0425_)
  );
  sky130_fd_sc_hd__or3_2 _2733_ (
    .A(_0396_),
    .B(_0146_),
    .C(_0141_),
    .X(_0426_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2734_ (
    .A1(_0391_),
    .A2(_0226_),
    .B1(_0424_),
    .C1(_0425_),
    .D1(_0426_),
    .Y(_0427_)
  );
  sky130_fd_sc_hd__or3_2 _2735_ (
    .A(_0400_),
    .B(_0239_),
    .C(_0240_),
    .X(_0428_)
  );
  sky130_fd_sc_hd__or3_2 _2736_ (
    .A(_0402_),
    .B(_0242_),
    .C(_0166_),
    .X(_0429_)
  );
  sky130_fd_sc_hd__or3_2 _2737_ (
    .A(_0404_),
    .B(_0309_),
    .C(_0148_),
    .X(_0430_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2738_ (
    .A1(_0399_),
    .A2(_0237_),
    .B1(_0428_),
    .C1(_0429_),
    .D1(_0430_),
    .Y(_0431_)
  );
  sky130_fd_sc_hd__or4_2 _2739_ (
    .A(_0421_),
    .B(_0423_),
    .C(_0427_),
    .D(_0431_),
    .X(_0432_)
  );
  sky130_fd_sc_hd__or4_2 _2740_ (
    .A(_0410_),
    .B(_0412_),
    .C(_0417_),
    .D(_0432_),
    .X(_0433_)
  );
  sky130_fd_sc_hd__buf_1 _2741_ (
    .A(_0433_),
    .X(\g_bit[2].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _2742_ (
    .A1(\g_bit[3].g_word[30].r_bit.Q ),
    .A2(_0023_),
    .A3(_0025_),
    .B1(_0030_),
    .B2(\g_bit[3].g_word[28].r_bit.Q ),
    .X(_0434_)
  );
  sky130_fd_sc_hd__a221o_2 _2743_ (
    .A1(\g_bit[3].g_word[4].r_bit.Q ),
    .A2(_0014_),
    .B1(_0021_),
    .B2(\g_bit[3].g_word[26].r_bit.Q ),
    .C1(_0434_),
    .X(_0435_)
  );
  sky130_fd_sc_hd__a22o_2 _2744_ (
    .A1(\g_bit[3].g_word[5].r_bit.Q ),
    .A2(_0043_),
    .B1(_0050_),
    .B2(\g_bit[3].g_word[2].r_bit.Q ),
    .X(_0436_)
  );
  sky130_fd_sc_hd__a221o_2 _2745_ (
    .A1(\g_bit[3].g_word[25].r_bit.Q ),
    .A2(_0035_),
    .B1(_0039_),
    .B2(\g_bit[3].g_word[31].r_bit.Q ),
    .C1(_0436_),
    .X(_0437_)
  );
  sky130_fd_sc_hd__a22o_2 _2746_ (
    .A1(\g_bit[3].g_word[13].r_bit.Q ),
    .A2(_0054_),
    .B1(_0057_),
    .B2(\g_bit[3].g_word[15].r_bit.Q ),
    .X(_0438_)
  );
  sky130_fd_sc_hd__a22o_2 _2747_ (
    .A1(\g_bit[3].g_word[11].r_bit.Q ),
    .A2(_0060_),
    .B1(_0062_),
    .B2(\g_bit[3].g_word[20].r_bit.Q ),
    .X(_0439_)
  );
  sky130_fd_sc_hd__a22o_2 _2748_ (
    .A1(\g_bit[3].g_word[19].r_bit.Q ),
    .A2(_0065_),
    .B1(_0067_),
    .B2(\g_bit[3].g_word[21].r_bit.Q ),
    .X(_0440_)
  );
  sky130_fd_sc_hd__a22o_2 _2749_ (
    .A1(\g_bit[3].g_word[17].r_bit.Q ),
    .A2(_0070_),
    .B1(_0072_),
    .B2(\g_bit[3].g_word[12].r_bit.Q ),
    .X(_0441_)
  );
  sky130_fd_sc_hd__or4_2 _2750_ (
    .A(_0438_),
    .B(_0439_),
    .C(_0440_),
    .D(_0441_),
    .X(_0442_)
  );
  sky130_fd_sc_hd__inv_2 _2751_ (
    .A(\g_bit[3].g_word[7].r_bit.Q ),
    .Y(_0443_)
  );
  sky130_fd_sc_hd__nor3_2 _2752_ (
    .A(_0443_),
    .B(_0082_),
    .C(_0004_),
    .Y(_0444_)
  );
  sky130_fd_sc_hd__inv_2 _2753_ (
    .A(\g_bit[3].g_word[3].r_bit.Q ),
    .Y(_0445_)
  );
  sky130_fd_sc_hd__nor3_2 _2754_ (
    .A(_0445_),
    .B(_0085_),
    .C(_0086_),
    .Y(_0446_)
  );
  sky130_fd_sc_hd__and3_2 _2755_ (
    .A(\g_bit[3].g_word[24].r_bit.Q ),
    .B(_0260_),
    .C(_0261_),
    .X(_0447_)
  );
  sky130_fd_sc_hd__a2111o_2 _2756_ (
    .A1(\g_bit[3].g_word[29].r_bit.Q ),
    .A2(_0076_),
    .B1(_0444_),
    .C1(_0446_),
    .D1(_0447_),
    .X(_0448_)
  );
  sky130_fd_sc_hd__and3_2 _2757_ (
    .A(\g_bit[3].g_word[27].r_bit.Q ),
    .B(_0094_),
    .C(_0095_),
    .X(_0449_)
  );
  sky130_fd_sc_hd__a221o_2 _2758_ (
    .A1(\g_bit[3].g_word[6].r_bit.Q ),
    .A2(_0090_),
    .B1(_0092_),
    .B2(\g_bit[3].g_word[1].r_bit.Q ),
    .C1(_0449_),
    .X(_0450_)
  );
  sky130_fd_sc_hd__inv_2 _2759_ (
    .A(\g_bit[3].g_word[23].r_bit.Q ),
    .Y(_0451_)
  );
  sky130_fd_sc_hd__inv_2 _2760_ (
    .A(\g_bit[3].g_word[10].r_bit.Q ),
    .Y(_0452_)
  );
  sky130_fd_sc_hd__buf_1 _2761_ (
    .A(_0015_),
    .X(_0453_)
  );
  sky130_fd_sc_hd__or3_2 _2762_ (
    .A(_0452_),
    .B(_0453_),
    .C(_0107_),
    .X(_0454_)
  );
  sky130_fd_sc_hd__inv_2 _2763_ (
    .A(\g_bit[3].g_word[9].r_bit.Q ),
    .Y(_0455_)
  );
  sky130_fd_sc_hd__or3_2 _2764_ (
    .A(_0455_),
    .B(_0106_),
    .C(_0110_),
    .X(_0456_)
  );
  sky130_fd_sc_hd__inv_2 _2765_ (
    .A(\g_bit[3].g_word[8].r_bit.Q ),
    .Y(_0457_)
  );
  sky130_fd_sc_hd__or3_2 _2766_ (
    .A(_0457_),
    .B(_0017_),
    .C(_0012_),
    .X(_0458_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2767_ (
    .A1(_0451_),
    .A2(_0101_),
    .B1(_0454_),
    .C1(_0456_),
    .D1(_0458_),
    .Y(_0459_)
  );
  sky130_fd_sc_hd__inv_2 _2768_ (
    .A(\g_bit[3].g_word[22].r_bit.Q ),
    .Y(_0460_)
  );
  sky130_fd_sc_hd__inv_2 _2769_ (
    .A(\g_bit[3].g_word[16].r_bit.Q ),
    .Y(_0461_)
  );
  sky130_fd_sc_hd__or3_2 _2770_ (
    .A(_0461_),
    .B(_0118_),
    .C(_0121_),
    .X(_0462_)
  );
  sky130_fd_sc_hd__inv_2 _2771_ (
    .A(\g_bit[3].g_word[14].r_bit.Q ),
    .Y(_0463_)
  );
  sky130_fd_sc_hd__or3_2 _2772_ (
    .A(_0463_),
    .B(_0124_),
    .C(_0037_),
    .X(_0464_)
  );
  sky130_fd_sc_hd__inv_2 _2773_ (
    .A(\g_bit[3].g_word[18].r_bit.Q ),
    .Y(_0465_)
  );
  sky130_fd_sc_hd__or3_2 _2774_ (
    .A(_0465_),
    .B(_0280_),
    .C(_0019_),
    .X(_0466_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2775_ (
    .A1(_0460_),
    .A2(_0116_),
    .B1(_0462_),
    .C1(_0464_),
    .D1(_0466_),
    .Y(_0467_)
  );
  sky130_fd_sc_hd__or4_2 _2776_ (
    .A(_0448_),
    .B(_0450_),
    .C(_0459_),
    .D(_0467_),
    .X(_0468_)
  );
  sky130_fd_sc_hd__or4_2 _2777_ (
    .A(_0435_),
    .B(_0437_),
    .C(_0442_),
    .D(_0468_),
    .X(_0469_)
  );
  sky130_fd_sc_hd__buf_1 _2778_ (
    .A(_0469_),
    .X(\g_bit[3].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _2779_ (
    .A1(\g_bit[3].g_word[30].r_bit.Q ),
    .A2(_0152_),
    .A3(_0154_),
    .B1(_0159_),
    .B2(\g_bit[3].g_word[28].r_bit.Q ),
    .X(_0470_)
  );
  sky130_fd_sc_hd__a221o_2 _2780_ (
    .A1(\g_bit[3].g_word[4].r_bit.Q ),
    .A2(_0143_),
    .B1(_0150_),
    .B2(\g_bit[3].g_word[26].r_bit.Q ),
    .C1(_0470_),
    .X(_0471_)
  );
  sky130_fd_sc_hd__a22o_2 _2781_ (
    .A1(\g_bit[3].g_word[5].r_bit.Q ),
    .A2(_0172_),
    .B1(_0179_),
    .B2(\g_bit[3].g_word[2].r_bit.Q ),
    .X(_0472_)
  );
  sky130_fd_sc_hd__a221o_2 _2782_ (
    .A1(\g_bit[3].g_word[25].r_bit.Q ),
    .A2(_0164_),
    .B1(_0168_),
    .B2(\g_bit[3].g_word[31].r_bit.Q ),
    .C1(_0472_),
    .X(_0473_)
  );
  sky130_fd_sc_hd__a22o_2 _2783_ (
    .A1(\g_bit[3].g_word[13].r_bit.Q ),
    .A2(_0183_),
    .B1(_0186_),
    .B2(\g_bit[3].g_word[15].r_bit.Q ),
    .X(_0474_)
  );
  sky130_fd_sc_hd__a22o_2 _2784_ (
    .A1(\g_bit[3].g_word[20].r_bit.Q ),
    .A2(_0189_),
    .B1(_0191_),
    .B2(\g_bit[3].g_word[11].r_bit.Q ),
    .X(_0475_)
  );
  sky130_fd_sc_hd__a22o_2 _2785_ (
    .A1(\g_bit[3].g_word[19].r_bit.Q ),
    .A2(_0194_),
    .B1(_0196_),
    .B2(\g_bit[3].g_word[21].r_bit.Q ),
    .X(_0476_)
  );
  sky130_fd_sc_hd__a22o_2 _2786_ (
    .A1(\g_bit[3].g_word[17].r_bit.Q ),
    .A2(_0199_),
    .B1(_0201_),
    .B2(\g_bit[3].g_word[12].r_bit.Q ),
    .X(_0477_)
  );
  sky130_fd_sc_hd__or4_2 _2787_ (
    .A(_0474_),
    .B(_0475_),
    .C(_0476_),
    .D(_0477_),
    .X(_0478_)
  );
  sky130_fd_sc_hd__nor3_2 _2788_ (
    .A(_0443_),
    .B(_0133_),
    .C(_0294_),
    .Y(_0479_)
  );
  sky130_fd_sc_hd__nor3_2 _2789_ (
    .A(_0445_),
    .B(_0212_),
    .C(_0210_),
    .Y(_0480_)
  );
  sky130_fd_sc_hd__and3_2 _2790_ (
    .A(\g_bit[3].g_word[24].r_bit.Q ),
    .B(_0297_),
    .C(_0298_),
    .X(_0481_)
  );
  sky130_fd_sc_hd__a2111o_2 _2791_ (
    .A1(\g_bit[3].g_word[29].r_bit.Q ),
    .A2(_0205_),
    .B1(_0479_),
    .C1(_0480_),
    .D1(_0481_),
    .X(_0482_)
  );
  sky130_fd_sc_hd__and3_2 _2792_ (
    .A(\g_bit[3].g_word[27].r_bit.Q ),
    .B(_0220_),
    .C(_0221_),
    .X(_0483_)
  );
  sky130_fd_sc_hd__a221o_2 _2793_ (
    .A1(\g_bit[3].g_word[6].r_bit.Q ),
    .A2(_0216_),
    .B1(_0218_),
    .B2(\g_bit[3].g_word[1].r_bit.Q ),
    .C1(_0483_),
    .X(_0484_)
  );
  sky130_fd_sc_hd__buf_1 _2794_ (
    .A(_0144_),
    .X(_0485_)
  );
  sky130_fd_sc_hd__or3_2 _2795_ (
    .A(_0452_),
    .B(_0485_),
    .C(_0230_),
    .X(_0486_)
  );
  sky130_fd_sc_hd__or3_2 _2796_ (
    .A(_0455_),
    .B(_0229_),
    .C(_0232_),
    .X(_0487_)
  );
  sky130_fd_sc_hd__or3_2 _2797_ (
    .A(_0457_),
    .B(_0146_),
    .C(_0141_),
    .X(_0488_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2798_ (
    .A1(_0451_),
    .A2(_0226_),
    .B1(_0486_),
    .C1(_0487_),
    .D1(_0488_),
    .Y(_0489_)
  );
  sky130_fd_sc_hd__or3_2 _2799_ (
    .A(_0461_),
    .B(_0239_),
    .C(_0240_),
    .X(_0490_)
  );
  sky130_fd_sc_hd__or3_2 _2800_ (
    .A(_0463_),
    .B(_0242_),
    .C(_0166_),
    .X(_0491_)
  );
  sky130_fd_sc_hd__or3_2 _2801_ (
    .A(_0465_),
    .B(_0309_),
    .C(_0148_),
    .X(_0492_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2802_ (
    .A1(_0460_),
    .A2(_0237_),
    .B1(_0490_),
    .C1(_0491_),
    .D1(_0492_),
    .Y(_0493_)
  );
  sky130_fd_sc_hd__or4_2 _2803_ (
    .A(_0482_),
    .B(_0484_),
    .C(_0489_),
    .D(_0493_),
    .X(_0494_)
  );
  sky130_fd_sc_hd__or4_2 _2804_ (
    .A(_0471_),
    .B(_0473_),
    .C(_0478_),
    .D(_0494_),
    .X(_0495_)
  );
  sky130_fd_sc_hd__buf_1 _2805_ (
    .A(_0495_),
    .X(\g_bit[3].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _2806_ (
    .A1(\g_bit[4].g_word[30].r_bit.Q ),
    .A2(_0023_),
    .A3(_0025_),
    .B1(_0030_),
    .B2(\g_bit[4].g_word[28].r_bit.Q ),
    .X(_0496_)
  );
  sky130_fd_sc_hd__a221o_2 _2807_ (
    .A1(\g_bit[4].g_word[4].r_bit.Q ),
    .A2(_0014_),
    .B1(_0021_),
    .B2(\g_bit[4].g_word[26].r_bit.Q ),
    .C1(_0496_),
    .X(_0497_)
  );
  sky130_fd_sc_hd__a22o_2 _2808_ (
    .A1(\g_bit[4].g_word[5].r_bit.Q ),
    .A2(_0043_),
    .B1(_0050_),
    .B2(\g_bit[4].g_word[2].r_bit.Q ),
    .X(_0498_)
  );
  sky130_fd_sc_hd__a221o_2 _2809_ (
    .A1(\g_bit[4].g_word[25].r_bit.Q ),
    .A2(_0035_),
    .B1(_0039_),
    .B2(\g_bit[4].g_word[31].r_bit.Q ),
    .C1(_0498_),
    .X(_0499_)
  );
  sky130_fd_sc_hd__a22o_2 _2810_ (
    .A1(\g_bit[4].g_word[13].r_bit.Q ),
    .A2(_0054_),
    .B1(_0057_),
    .B2(\g_bit[4].g_word[15].r_bit.Q ),
    .X(_0500_)
  );
  sky130_fd_sc_hd__a22o_2 _2811_ (
    .A1(\g_bit[4].g_word[11].r_bit.Q ),
    .A2(_0060_),
    .B1(_0062_),
    .B2(\g_bit[4].g_word[20].r_bit.Q ),
    .X(_0501_)
  );
  sky130_fd_sc_hd__a22o_2 _2812_ (
    .A1(\g_bit[4].g_word[19].r_bit.Q ),
    .A2(_0065_),
    .B1(_0067_),
    .B2(\g_bit[4].g_word[21].r_bit.Q ),
    .X(_0502_)
  );
  sky130_fd_sc_hd__a22o_2 _2813_ (
    .A1(\g_bit[4].g_word[17].r_bit.Q ),
    .A2(_0070_),
    .B1(_0072_),
    .B2(\g_bit[4].g_word[12].r_bit.Q ),
    .X(_0503_)
  );
  sky130_fd_sc_hd__or4_2 _2814_ (
    .A(_0500_),
    .B(_0501_),
    .C(_0502_),
    .D(_0503_),
    .X(_0504_)
  );
  sky130_fd_sc_hd__inv_2 _2815_ (
    .A(\g_bit[4].g_word[7].r_bit.Q ),
    .Y(_0505_)
  );
  sky130_fd_sc_hd__nor3_2 _2816_ (
    .A(_0505_),
    .B(_0082_),
    .C(_0004_),
    .Y(_0506_)
  );
  sky130_fd_sc_hd__inv_2 _2817_ (
    .A(\g_bit[4].g_word[3].r_bit.Q ),
    .Y(_0507_)
  );
  sky130_fd_sc_hd__nor3_2 _2818_ (
    .A(_0507_),
    .B(_0085_),
    .C(_0086_),
    .Y(_0508_)
  );
  sky130_fd_sc_hd__and3_2 _2819_ (
    .A(\g_bit[4].g_word[24].r_bit.Q ),
    .B(_0260_),
    .C(_0261_),
    .X(_0509_)
  );
  sky130_fd_sc_hd__a2111o_2 _2820_ (
    .A1(\g_bit[4].g_word[29].r_bit.Q ),
    .A2(_0076_),
    .B1(_0506_),
    .C1(_0508_),
    .D1(_0509_),
    .X(_0510_)
  );
  sky130_fd_sc_hd__and3_2 _2821_ (
    .A(\g_bit[4].g_word[27].r_bit.Q ),
    .B(_0094_),
    .C(_0095_),
    .X(_0511_)
  );
  sky130_fd_sc_hd__a221o_2 _2822_ (
    .A1(\g_bit[4].g_word[6].r_bit.Q ),
    .A2(_0090_),
    .B1(_0092_),
    .B2(\g_bit[4].g_word[1].r_bit.Q ),
    .C1(_0511_),
    .X(_0512_)
  );
  sky130_fd_sc_hd__inv_2 _2823_ (
    .A(\g_bit[4].g_word[23].r_bit.Q ),
    .Y(_0513_)
  );
  sky130_fd_sc_hd__inv_2 _2824_ (
    .A(\g_bit[4].g_word[10].r_bit.Q ),
    .Y(_0514_)
  );
  sky130_fd_sc_hd__or3_2 _2825_ (
    .A(_0514_),
    .B(_0453_),
    .C(_0107_),
    .X(_0515_)
  );
  sky130_fd_sc_hd__inv_2 _2826_ (
    .A(\g_bit[4].g_word[9].r_bit.Q ),
    .Y(_0516_)
  );
  sky130_fd_sc_hd__or3_2 _2827_ (
    .A(_0516_),
    .B(_0106_),
    .C(_0110_),
    .X(_0517_)
  );
  sky130_fd_sc_hd__inv_2 _2828_ (
    .A(\g_bit[4].g_word[8].r_bit.Q ),
    .Y(_0518_)
  );
  sky130_fd_sc_hd__or3_2 _2829_ (
    .A(_0518_),
    .B(_0017_),
    .C(_0012_),
    .X(_0519_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2830_ (
    .A1(_0513_),
    .A2(_0101_),
    .B1(_0515_),
    .C1(_0517_),
    .D1(_0519_),
    .Y(_0520_)
  );
  sky130_fd_sc_hd__inv_2 _2831_ (
    .A(\g_bit[4].g_word[22].r_bit.Q ),
    .Y(_0521_)
  );
  sky130_fd_sc_hd__inv_2 _2832_ (
    .A(\g_bit[4].g_word[16].r_bit.Q ),
    .Y(_0522_)
  );
  sky130_fd_sc_hd__or3_2 _2833_ (
    .A(_0522_),
    .B(_0118_),
    .C(_0121_),
    .X(_0523_)
  );
  sky130_fd_sc_hd__inv_2 _2834_ (
    .A(\g_bit[4].g_word[14].r_bit.Q ),
    .Y(_0524_)
  );
  sky130_fd_sc_hd__or3_2 _2835_ (
    .A(_0524_),
    .B(_0124_),
    .C(_0037_),
    .X(_0525_)
  );
  sky130_fd_sc_hd__inv_2 _2836_ (
    .A(\g_bit[4].g_word[18].r_bit.Q ),
    .Y(_0526_)
  );
  sky130_fd_sc_hd__or3_2 _2837_ (
    .A(_0526_),
    .B(_0280_),
    .C(_0019_),
    .X(_0527_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2838_ (
    .A1(_0521_),
    .A2(_0116_),
    .B1(_0523_),
    .C1(_0525_),
    .D1(_0527_),
    .Y(_0528_)
  );
  sky130_fd_sc_hd__or4_2 _2839_ (
    .A(_0510_),
    .B(_0512_),
    .C(_0520_),
    .D(_0528_),
    .X(_0529_)
  );
  sky130_fd_sc_hd__or4_2 _2840_ (
    .A(_0497_),
    .B(_0499_),
    .C(_0504_),
    .D(_0529_),
    .X(_0530_)
  );
  sky130_fd_sc_hd__buf_1 _2841_ (
    .A(_0530_),
    .X(\g_bit[4].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _2842_ (
    .A1(\g_bit[4].g_word[30].r_bit.Q ),
    .A2(_0152_),
    .A3(_0154_),
    .B1(_0159_),
    .B2(\g_bit[4].g_word[28].r_bit.Q ),
    .X(_0531_)
  );
  sky130_fd_sc_hd__a221o_2 _2843_ (
    .A1(\g_bit[4].g_word[4].r_bit.Q ),
    .A2(_0143_),
    .B1(_0150_),
    .B2(\g_bit[4].g_word[26].r_bit.Q ),
    .C1(_0531_),
    .X(_0532_)
  );
  sky130_fd_sc_hd__a22o_2 _2844_ (
    .A1(\g_bit[4].g_word[5].r_bit.Q ),
    .A2(_0172_),
    .B1(_0179_),
    .B2(\g_bit[4].g_word[2].r_bit.Q ),
    .X(_0533_)
  );
  sky130_fd_sc_hd__a221o_2 _2845_ (
    .A1(\g_bit[4].g_word[25].r_bit.Q ),
    .A2(_0164_),
    .B1(_0168_),
    .B2(\g_bit[4].g_word[31].r_bit.Q ),
    .C1(_0533_),
    .X(_0534_)
  );
  sky130_fd_sc_hd__a22o_2 _2846_ (
    .A1(\g_bit[4].g_word[13].r_bit.Q ),
    .A2(_0183_),
    .B1(_0186_),
    .B2(\g_bit[4].g_word[15].r_bit.Q ),
    .X(_0535_)
  );
  sky130_fd_sc_hd__a22o_2 _2847_ (
    .A1(\g_bit[4].g_word[20].r_bit.Q ),
    .A2(_0189_),
    .B1(_0191_),
    .B2(\g_bit[4].g_word[11].r_bit.Q ),
    .X(_0536_)
  );
  sky130_fd_sc_hd__a22o_2 _2848_ (
    .A1(\g_bit[4].g_word[19].r_bit.Q ),
    .A2(_0194_),
    .B1(_0196_),
    .B2(\g_bit[4].g_word[21].r_bit.Q ),
    .X(_0537_)
  );
  sky130_fd_sc_hd__a22o_2 _2849_ (
    .A1(\g_bit[4].g_word[17].r_bit.Q ),
    .A2(_0199_),
    .B1(_0201_),
    .B2(\g_bit[4].g_word[12].r_bit.Q ),
    .X(_0538_)
  );
  sky130_fd_sc_hd__or4_2 _2850_ (
    .A(_0535_),
    .B(_0536_),
    .C(_0537_),
    .D(_0538_),
    .X(_0539_)
  );
  sky130_fd_sc_hd__nor3_2 _2851_ (
    .A(_0505_),
    .B(_0133_),
    .C(_0294_),
    .Y(_0540_)
  );
  sky130_fd_sc_hd__nor3_2 _2852_ (
    .A(_0507_),
    .B(_0212_),
    .C(_0210_),
    .Y(_0541_)
  );
  sky130_fd_sc_hd__and3_2 _2853_ (
    .A(\g_bit[4].g_word[24].r_bit.Q ),
    .B(_0297_),
    .C(_0298_),
    .X(_0542_)
  );
  sky130_fd_sc_hd__a2111o_2 _2854_ (
    .A1(\g_bit[4].g_word[29].r_bit.Q ),
    .A2(_0205_),
    .B1(_0540_),
    .C1(_0541_),
    .D1(_0542_),
    .X(_0543_)
  );
  sky130_fd_sc_hd__and3_2 _2855_ (
    .A(\g_bit[4].g_word[27].r_bit.Q ),
    .B(_0220_),
    .C(_0221_),
    .X(_0544_)
  );
  sky130_fd_sc_hd__a221o_2 _2856_ (
    .A1(\g_bit[4].g_word[6].r_bit.Q ),
    .A2(_0216_),
    .B1(_0218_),
    .B2(\g_bit[4].g_word[1].r_bit.Q ),
    .C1(_0544_),
    .X(_0545_)
  );
  sky130_fd_sc_hd__or3_2 _2857_ (
    .A(_0514_),
    .B(_0485_),
    .C(_0230_),
    .X(_0546_)
  );
  sky130_fd_sc_hd__or3_2 _2858_ (
    .A(_0516_),
    .B(_0229_),
    .C(_0232_),
    .X(_0547_)
  );
  sky130_fd_sc_hd__or3_2 _2859_ (
    .A(_0518_),
    .B(_0146_),
    .C(_0141_),
    .X(_0548_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2860_ (
    .A1(_0513_),
    .A2(_0226_),
    .B1(_0546_),
    .C1(_0547_),
    .D1(_0548_),
    .Y(_0549_)
  );
  sky130_fd_sc_hd__or3_2 _2861_ (
    .A(_0522_),
    .B(_0239_),
    .C(_0240_),
    .X(_0550_)
  );
  sky130_fd_sc_hd__or3_2 _2862_ (
    .A(_0524_),
    .B(_0242_),
    .C(_0166_),
    .X(_0551_)
  );
  sky130_fd_sc_hd__or3_2 _2863_ (
    .A(_0526_),
    .B(_0309_),
    .C(_0148_),
    .X(_0552_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2864_ (
    .A1(_0521_),
    .A2(_0237_),
    .B1(_0550_),
    .C1(_0551_),
    .D1(_0552_),
    .Y(_0553_)
  );
  sky130_fd_sc_hd__or4_2 _2865_ (
    .A(_0543_),
    .B(_0545_),
    .C(_0549_),
    .D(_0553_),
    .X(_0554_)
  );
  sky130_fd_sc_hd__or4_2 _2866_ (
    .A(_0532_),
    .B(_0534_),
    .C(_0539_),
    .D(_0554_),
    .X(_0555_)
  );
  sky130_fd_sc_hd__buf_1 _2867_ (
    .A(_0555_),
    .X(\g_bit[4].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _2868_ (
    .A1(\g_bit[5].g_word[30].r_bit.Q ),
    .A2(_0023_),
    .A3(_0025_),
    .B1(_0030_),
    .B2(\g_bit[5].g_word[28].r_bit.Q ),
    .X(_0556_)
  );
  sky130_fd_sc_hd__a221o_2 _2869_ (
    .A1(\g_bit[5].g_word[4].r_bit.Q ),
    .A2(_0014_),
    .B1(_0021_),
    .B2(\g_bit[5].g_word[26].r_bit.Q ),
    .C1(_0556_),
    .X(_0557_)
  );
  sky130_fd_sc_hd__a22o_2 _2870_ (
    .A1(\g_bit[5].g_word[5].r_bit.Q ),
    .A2(_0043_),
    .B1(_0050_),
    .B2(\g_bit[5].g_word[2].r_bit.Q ),
    .X(_0558_)
  );
  sky130_fd_sc_hd__a221o_2 _2871_ (
    .A1(\g_bit[5].g_word[25].r_bit.Q ),
    .A2(_0035_),
    .B1(_0039_),
    .B2(\g_bit[5].g_word[31].r_bit.Q ),
    .C1(_0558_),
    .X(_0559_)
  );
  sky130_fd_sc_hd__a22o_2 _2872_ (
    .A1(\g_bit[5].g_word[13].r_bit.Q ),
    .A2(_0054_),
    .B1(_0057_),
    .B2(\g_bit[5].g_word[15].r_bit.Q ),
    .X(_0560_)
  );
  sky130_fd_sc_hd__a22o_2 _2873_ (
    .A1(\g_bit[5].g_word[11].r_bit.Q ),
    .A2(_0060_),
    .B1(_0062_),
    .B2(\g_bit[5].g_word[20].r_bit.Q ),
    .X(_0561_)
  );
  sky130_fd_sc_hd__a22o_2 _2874_ (
    .A1(\g_bit[5].g_word[19].r_bit.Q ),
    .A2(_0065_),
    .B1(_0067_),
    .B2(\g_bit[5].g_word[21].r_bit.Q ),
    .X(_0562_)
  );
  sky130_fd_sc_hd__a22o_2 _2875_ (
    .A1(\g_bit[5].g_word[17].r_bit.Q ),
    .A2(_0070_),
    .B1(_0072_),
    .B2(\g_bit[5].g_word[12].r_bit.Q ),
    .X(_0563_)
  );
  sky130_fd_sc_hd__or4_2 _2876_ (
    .A(_0560_),
    .B(_0561_),
    .C(_0562_),
    .D(_0563_),
    .X(_0564_)
  );
  sky130_fd_sc_hd__inv_2 _2877_ (
    .A(\g_bit[5].g_word[7].r_bit.Q ),
    .Y(_0565_)
  );
  sky130_fd_sc_hd__nor3_2 _2878_ (
    .A(_0565_),
    .B(_0082_),
    .C(_0004_),
    .Y(_0566_)
  );
  sky130_fd_sc_hd__inv_2 _2879_ (
    .A(\g_bit[5].g_word[3].r_bit.Q ),
    .Y(_0567_)
  );
  sky130_fd_sc_hd__nor3_2 _2880_ (
    .A(_0567_),
    .B(_0085_),
    .C(_0086_),
    .Y(_0568_)
  );
  sky130_fd_sc_hd__and3_2 _2881_ (
    .A(\g_bit[5].g_word[24].r_bit.Q ),
    .B(_0260_),
    .C(_0261_),
    .X(_0569_)
  );
  sky130_fd_sc_hd__a2111o_2 _2882_ (
    .A1(\g_bit[5].g_word[29].r_bit.Q ),
    .A2(_0076_),
    .B1(_0566_),
    .C1(_0568_),
    .D1(_0569_),
    .X(_0570_)
  );
  sky130_fd_sc_hd__and3_2 _2883_ (
    .A(\g_bit[5].g_word[27].r_bit.Q ),
    .B(_0094_),
    .C(_0095_),
    .X(_0571_)
  );
  sky130_fd_sc_hd__a221o_2 _2884_ (
    .A1(\g_bit[5].g_word[6].r_bit.Q ),
    .A2(_0090_),
    .B1(_0092_),
    .B2(\g_bit[5].g_word[1].r_bit.Q ),
    .C1(_0571_),
    .X(_0572_)
  );
  sky130_fd_sc_hd__inv_2 _2885_ (
    .A(\g_bit[5].g_word[23].r_bit.Q ),
    .Y(_0573_)
  );
  sky130_fd_sc_hd__inv_2 _2886_ (
    .A(\g_bit[5].g_word[10].r_bit.Q ),
    .Y(_0574_)
  );
  sky130_fd_sc_hd__or3_2 _2887_ (
    .A(_0574_),
    .B(_0453_),
    .C(_0107_),
    .X(_0575_)
  );
  sky130_fd_sc_hd__inv_2 _2888_ (
    .A(\g_bit[5].g_word[9].r_bit.Q ),
    .Y(_0576_)
  );
  sky130_fd_sc_hd__buf_1 _2889_ (
    .A(_0015_),
    .X(_0577_)
  );
  sky130_fd_sc_hd__or3_2 _2890_ (
    .A(_0576_),
    .B(_0577_),
    .C(_0110_),
    .X(_0578_)
  );
  sky130_fd_sc_hd__inv_2 _2891_ (
    .A(\g_bit[5].g_word[8].r_bit.Q ),
    .Y(_0579_)
  );
  sky130_fd_sc_hd__or3_2 _2892_ (
    .A(_0579_),
    .B(_0017_),
    .C(_0012_),
    .X(_0580_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2893_ (
    .A1(_0573_),
    .A2(_0101_),
    .B1(_0575_),
    .C1(_0578_),
    .D1(_0580_),
    .Y(_0581_)
  );
  sky130_fd_sc_hd__inv_2 _2894_ (
    .A(\g_bit[5].g_word[22].r_bit.Q ),
    .Y(_0582_)
  );
  sky130_fd_sc_hd__inv_2 _2895_ (
    .A(\g_bit[5].g_word[16].r_bit.Q ),
    .Y(_0583_)
  );
  sky130_fd_sc_hd__buf_1 _2896_ (
    .A(_0045_),
    .X(_0584_)
  );
  sky130_fd_sc_hd__or3_2 _2897_ (
    .A(_0583_),
    .B(_0584_),
    .C(_0121_),
    .X(_0585_)
  );
  sky130_fd_sc_hd__inv_2 _2898_ (
    .A(\g_bit[5].g_word[14].r_bit.Q ),
    .Y(_0586_)
  );
  sky130_fd_sc_hd__or3_2 _2899_ (
    .A(_0586_),
    .B(_0124_),
    .C(_0037_),
    .X(_0587_)
  );
  sky130_fd_sc_hd__inv_2 _2900_ (
    .A(\g_bit[5].g_word[18].r_bit.Q ),
    .Y(_0588_)
  );
  sky130_fd_sc_hd__or3_2 _2901_ (
    .A(_0588_),
    .B(_0280_),
    .C(_0019_),
    .X(_0589_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2902_ (
    .A1(_0582_),
    .A2(_0116_),
    .B1(_0585_),
    .C1(_0587_),
    .D1(_0589_),
    .Y(_0590_)
  );
  sky130_fd_sc_hd__or4_2 _2903_ (
    .A(_0570_),
    .B(_0572_),
    .C(_0581_),
    .D(_0590_),
    .X(_0591_)
  );
  sky130_fd_sc_hd__or4_2 _2904_ (
    .A(_0557_),
    .B(_0559_),
    .C(_0564_),
    .D(_0591_),
    .X(_0592_)
  );
  sky130_fd_sc_hd__buf_1 _2905_ (
    .A(_0592_),
    .X(\g_bit[5].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _2906_ (
    .A1(\g_bit[5].g_word[30].r_bit.Q ),
    .A2(_0152_),
    .A3(_0154_),
    .B1(_0159_),
    .B2(\g_bit[5].g_word[28].r_bit.Q ),
    .X(_0593_)
  );
  sky130_fd_sc_hd__a221o_2 _2907_ (
    .A1(\g_bit[5].g_word[4].r_bit.Q ),
    .A2(_0143_),
    .B1(_0150_),
    .B2(\g_bit[5].g_word[26].r_bit.Q ),
    .C1(_0593_),
    .X(_0594_)
  );
  sky130_fd_sc_hd__a22o_2 _2908_ (
    .A1(\g_bit[5].g_word[5].r_bit.Q ),
    .A2(_0172_),
    .B1(_0179_),
    .B2(\g_bit[5].g_word[2].r_bit.Q ),
    .X(_0595_)
  );
  sky130_fd_sc_hd__a221o_2 _2909_ (
    .A1(\g_bit[5].g_word[25].r_bit.Q ),
    .A2(_0164_),
    .B1(_0168_),
    .B2(\g_bit[5].g_word[31].r_bit.Q ),
    .C1(_0595_),
    .X(_0596_)
  );
  sky130_fd_sc_hd__a22o_2 _2910_ (
    .A1(\g_bit[5].g_word[13].r_bit.Q ),
    .A2(_0183_),
    .B1(_0186_),
    .B2(\g_bit[5].g_word[15].r_bit.Q ),
    .X(_0597_)
  );
  sky130_fd_sc_hd__a22o_2 _2911_ (
    .A1(\g_bit[5].g_word[20].r_bit.Q ),
    .A2(_0189_),
    .B1(_0191_),
    .B2(\g_bit[5].g_word[11].r_bit.Q ),
    .X(_0598_)
  );
  sky130_fd_sc_hd__a22o_2 _2912_ (
    .A1(\g_bit[5].g_word[19].r_bit.Q ),
    .A2(_0194_),
    .B1(_0196_),
    .B2(\g_bit[5].g_word[21].r_bit.Q ),
    .X(_0599_)
  );
  sky130_fd_sc_hd__a22o_2 _2913_ (
    .A1(\g_bit[5].g_word[17].r_bit.Q ),
    .A2(_0199_),
    .B1(_0201_),
    .B2(\g_bit[5].g_word[12].r_bit.Q ),
    .X(_0600_)
  );
  sky130_fd_sc_hd__or4_2 _2914_ (
    .A(_0597_),
    .B(_0598_),
    .C(_0599_),
    .D(_0600_),
    .X(_0601_)
  );
  sky130_fd_sc_hd__nor3_2 _2915_ (
    .A(_0565_),
    .B(_0133_),
    .C(_0294_),
    .Y(_0602_)
  );
  sky130_fd_sc_hd__nor3_2 _2916_ (
    .A(_0567_),
    .B(_0212_),
    .C(_0210_),
    .Y(_0603_)
  );
  sky130_fd_sc_hd__and3_2 _2917_ (
    .A(\g_bit[5].g_word[24].r_bit.Q ),
    .B(_0297_),
    .C(_0298_),
    .X(_0604_)
  );
  sky130_fd_sc_hd__a2111o_2 _2918_ (
    .A1(\g_bit[5].g_word[29].r_bit.Q ),
    .A2(_0205_),
    .B1(_0602_),
    .C1(_0603_),
    .D1(_0604_),
    .X(_0605_)
  );
  sky130_fd_sc_hd__and3_2 _2919_ (
    .A(\g_bit[5].g_word[27].r_bit.Q ),
    .B(_0220_),
    .C(_0221_),
    .X(_0606_)
  );
  sky130_fd_sc_hd__a221o_2 _2920_ (
    .A1(\g_bit[5].g_word[6].r_bit.Q ),
    .A2(_0216_),
    .B1(_0218_),
    .B2(\g_bit[5].g_word[1].r_bit.Q ),
    .C1(_0606_),
    .X(_0607_)
  );
  sky130_fd_sc_hd__or3_2 _2921_ (
    .A(_0574_),
    .B(_0485_),
    .C(_0230_),
    .X(_0608_)
  );
  sky130_fd_sc_hd__buf_1 _2922_ (
    .A(_0144_),
    .X(_0609_)
  );
  sky130_fd_sc_hd__or3_2 _2923_ (
    .A(_0576_),
    .B(_0609_),
    .C(_0232_),
    .X(_0610_)
  );
  sky130_fd_sc_hd__or3_2 _2924_ (
    .A(_0579_),
    .B(_0146_),
    .C(_0141_),
    .X(_0611_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2925_ (
    .A1(_0573_),
    .A2(_0226_),
    .B1(_0608_),
    .C1(_0610_),
    .D1(_0611_),
    .Y(_0612_)
  );
  sky130_fd_sc_hd__or3_2 _2926_ (
    .A(_0583_),
    .B(_0239_),
    .C(_0240_),
    .X(_0613_)
  );
  sky130_fd_sc_hd__or3_2 _2927_ (
    .A(_0586_),
    .B(_0242_),
    .C(_0166_),
    .X(_0614_)
  );
  sky130_fd_sc_hd__or3_2 _2928_ (
    .A(_0588_),
    .B(_0309_),
    .C(_0148_),
    .X(_0615_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2929_ (
    .A1(_0582_),
    .A2(_0237_),
    .B1(_0613_),
    .C1(_0614_),
    .D1(_0615_),
    .Y(_0616_)
  );
  sky130_fd_sc_hd__or4_2 _2930_ (
    .A(_0605_),
    .B(_0607_),
    .C(_0612_),
    .D(_0616_),
    .X(_0617_)
  );
  sky130_fd_sc_hd__or4_2 _2931_ (
    .A(_0594_),
    .B(_0596_),
    .C(_0601_),
    .D(_0617_),
    .X(_0618_)
  );
  sky130_fd_sc_hd__buf_1 _2932_ (
    .A(_0618_),
    .X(\g_bit[5].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _2933_ (
    .A1(\g_bit[6].g_word[30].r_bit.Q ),
    .A2(_0023_),
    .A3(_0025_),
    .B1(_0030_),
    .B2(\g_bit[6].g_word[28].r_bit.Q ),
    .X(_0619_)
  );
  sky130_fd_sc_hd__a221o_2 _2934_ (
    .A1(\g_bit[6].g_word[4].r_bit.Q ),
    .A2(_0014_),
    .B1(_0021_),
    .B2(\g_bit[6].g_word[26].r_bit.Q ),
    .C1(_0619_),
    .X(_0620_)
  );
  sky130_fd_sc_hd__a22o_2 _2935_ (
    .A1(\g_bit[6].g_word[5].r_bit.Q ),
    .A2(_0043_),
    .B1(_0050_),
    .B2(\g_bit[6].g_word[2].r_bit.Q ),
    .X(_0621_)
  );
  sky130_fd_sc_hd__a221o_2 _2936_ (
    .A1(\g_bit[6].g_word[25].r_bit.Q ),
    .A2(_0035_),
    .B1(_0039_),
    .B2(\g_bit[6].g_word[31].r_bit.Q ),
    .C1(_0621_),
    .X(_0622_)
  );
  sky130_fd_sc_hd__a22o_2 _2937_ (
    .A1(\g_bit[6].g_word[13].r_bit.Q ),
    .A2(_0054_),
    .B1(_0057_),
    .B2(\g_bit[6].g_word[15].r_bit.Q ),
    .X(_0623_)
  );
  sky130_fd_sc_hd__a22o_2 _2938_ (
    .A1(\g_bit[6].g_word[11].r_bit.Q ),
    .A2(_0060_),
    .B1(_0062_),
    .B2(\g_bit[6].g_word[20].r_bit.Q ),
    .X(_0624_)
  );
  sky130_fd_sc_hd__a22o_2 _2939_ (
    .A1(\g_bit[6].g_word[19].r_bit.Q ),
    .A2(_0065_),
    .B1(_0067_),
    .B2(\g_bit[6].g_word[21].r_bit.Q ),
    .X(_0625_)
  );
  sky130_fd_sc_hd__a22o_2 _2940_ (
    .A1(\g_bit[6].g_word[17].r_bit.Q ),
    .A2(_0070_),
    .B1(_0072_),
    .B2(\g_bit[6].g_word[12].r_bit.Q ),
    .X(_0626_)
  );
  sky130_fd_sc_hd__or4_2 _2941_ (
    .A(_0623_),
    .B(_0624_),
    .C(_0625_),
    .D(_0626_),
    .X(_0627_)
  );
  sky130_fd_sc_hd__inv_2 _2942_ (
    .A(\g_bit[6].g_word[7].r_bit.Q ),
    .Y(_0628_)
  );
  sky130_fd_sc_hd__nor3_2 _2943_ (
    .A(_0628_),
    .B(_0082_),
    .C(_0004_),
    .Y(_0629_)
  );
  sky130_fd_sc_hd__inv_2 _2944_ (
    .A(\g_bit[6].g_word[3].r_bit.Q ),
    .Y(_0630_)
  );
  sky130_fd_sc_hd__nor3_2 _2945_ (
    .A(_0630_),
    .B(_0085_),
    .C(_0086_),
    .Y(_0631_)
  );
  sky130_fd_sc_hd__and3_2 _2946_ (
    .A(\g_bit[6].g_word[24].r_bit.Q ),
    .B(_0260_),
    .C(_0261_),
    .X(_0632_)
  );
  sky130_fd_sc_hd__a2111o_2 _2947_ (
    .A1(\g_bit[6].g_word[29].r_bit.Q ),
    .A2(_0076_),
    .B1(_0629_),
    .C1(_0631_),
    .D1(_0632_),
    .X(_0633_)
  );
  sky130_fd_sc_hd__and3_2 _2948_ (
    .A(\g_bit[6].g_word[27].r_bit.Q ),
    .B(_0094_),
    .C(_0095_),
    .X(_0634_)
  );
  sky130_fd_sc_hd__a221o_2 _2949_ (
    .A1(\g_bit[6].g_word[6].r_bit.Q ),
    .A2(_0090_),
    .B1(_0092_),
    .B2(\g_bit[6].g_word[1].r_bit.Q ),
    .C1(_0634_),
    .X(_0635_)
  );
  sky130_fd_sc_hd__inv_2 _2950_ (
    .A(\g_bit[6].g_word[23].r_bit.Q ),
    .Y(_0636_)
  );
  sky130_fd_sc_hd__inv_2 _2951_ (
    .A(\g_bit[6].g_word[10].r_bit.Q ),
    .Y(_0637_)
  );
  sky130_fd_sc_hd__or3_2 _2952_ (
    .A(_0637_),
    .B(_0453_),
    .C(_0107_),
    .X(_0638_)
  );
  sky130_fd_sc_hd__inv_2 _2953_ (
    .A(\g_bit[6].g_word[9].r_bit.Q ),
    .Y(_0639_)
  );
  sky130_fd_sc_hd__or3_2 _2954_ (
    .A(_0639_),
    .B(_0577_),
    .C(_0110_),
    .X(_0640_)
  );
  sky130_fd_sc_hd__inv_2 _2955_ (
    .A(\g_bit[6].g_word[8].r_bit.Q ),
    .Y(_0641_)
  );
  sky130_fd_sc_hd__or3_2 _2956_ (
    .A(_0641_),
    .B(_0017_),
    .C(_0012_),
    .X(_0642_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2957_ (
    .A1(_0636_),
    .A2(_0101_),
    .B1(_0638_),
    .C1(_0640_),
    .D1(_0642_),
    .Y(_0643_)
  );
  sky130_fd_sc_hd__inv_2 _2958_ (
    .A(\g_bit[6].g_word[22].r_bit.Q ),
    .Y(_0644_)
  );
  sky130_fd_sc_hd__inv_2 _2959_ (
    .A(\g_bit[6].g_word[16].r_bit.Q ),
    .Y(_0645_)
  );
  sky130_fd_sc_hd__or3_2 _2960_ (
    .A(_0645_),
    .B(_0584_),
    .C(_0121_),
    .X(_0646_)
  );
  sky130_fd_sc_hd__inv_2 _2961_ (
    .A(\g_bit[6].g_word[14].r_bit.Q ),
    .Y(_0647_)
  );
  sky130_fd_sc_hd__or3_2 _2962_ (
    .A(_0647_),
    .B(_0124_),
    .C(_0037_),
    .X(_0648_)
  );
  sky130_fd_sc_hd__inv_2 _2963_ (
    .A(\g_bit[6].g_word[18].r_bit.Q ),
    .Y(_0649_)
  );
  sky130_fd_sc_hd__or3_2 _2964_ (
    .A(_0649_),
    .B(_0280_),
    .C(_0019_),
    .X(_0650_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2965_ (
    .A1(_0644_),
    .A2(_0116_),
    .B1(_0646_),
    .C1(_0648_),
    .D1(_0650_),
    .Y(_0651_)
  );
  sky130_fd_sc_hd__or4_2 _2966_ (
    .A(_0633_),
    .B(_0635_),
    .C(_0643_),
    .D(_0651_),
    .X(_0652_)
  );
  sky130_fd_sc_hd__or4_2 _2967_ (
    .A(_0620_),
    .B(_0622_),
    .C(_0627_),
    .D(_0652_),
    .X(_0653_)
  );
  sky130_fd_sc_hd__buf_1 _2968_ (
    .A(_0653_),
    .X(\g_bit[6].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _2969_ (
    .A1(\g_bit[6].g_word[30].r_bit.Q ),
    .A2(_0152_),
    .A3(_0154_),
    .B1(_0159_),
    .B2(\g_bit[6].g_word[28].r_bit.Q ),
    .X(_0654_)
  );
  sky130_fd_sc_hd__a221o_2 _2970_ (
    .A1(\g_bit[6].g_word[4].r_bit.Q ),
    .A2(_0143_),
    .B1(_0150_),
    .B2(\g_bit[6].g_word[26].r_bit.Q ),
    .C1(_0654_),
    .X(_0655_)
  );
  sky130_fd_sc_hd__a22o_2 _2971_ (
    .A1(\g_bit[6].g_word[5].r_bit.Q ),
    .A2(_0172_),
    .B1(_0179_),
    .B2(\g_bit[6].g_word[2].r_bit.Q ),
    .X(_0656_)
  );
  sky130_fd_sc_hd__a221o_2 _2972_ (
    .A1(\g_bit[6].g_word[25].r_bit.Q ),
    .A2(_0164_),
    .B1(_0168_),
    .B2(\g_bit[6].g_word[31].r_bit.Q ),
    .C1(_0656_),
    .X(_0657_)
  );
  sky130_fd_sc_hd__a22o_2 _2973_ (
    .A1(\g_bit[6].g_word[13].r_bit.Q ),
    .A2(_0183_),
    .B1(_0186_),
    .B2(\g_bit[6].g_word[15].r_bit.Q ),
    .X(_0658_)
  );
  sky130_fd_sc_hd__a22o_2 _2974_ (
    .A1(\g_bit[6].g_word[20].r_bit.Q ),
    .A2(_0189_),
    .B1(_0191_),
    .B2(\g_bit[6].g_word[11].r_bit.Q ),
    .X(_0659_)
  );
  sky130_fd_sc_hd__a22o_2 _2975_ (
    .A1(\g_bit[6].g_word[19].r_bit.Q ),
    .A2(_0194_),
    .B1(_0196_),
    .B2(\g_bit[6].g_word[21].r_bit.Q ),
    .X(_0660_)
  );
  sky130_fd_sc_hd__a22o_2 _2976_ (
    .A1(\g_bit[6].g_word[17].r_bit.Q ),
    .A2(_0199_),
    .B1(_0201_),
    .B2(\g_bit[6].g_word[12].r_bit.Q ),
    .X(_0661_)
  );
  sky130_fd_sc_hd__or4_2 _2977_ (
    .A(_0658_),
    .B(_0659_),
    .C(_0660_),
    .D(_0661_),
    .X(_0662_)
  );
  sky130_fd_sc_hd__nor3_2 _2978_ (
    .A(_0628_),
    .B(_0133_),
    .C(_0294_),
    .Y(_0663_)
  );
  sky130_fd_sc_hd__nor3_2 _2979_ (
    .A(_0630_),
    .B(_0212_),
    .C(_0210_),
    .Y(_0664_)
  );
  sky130_fd_sc_hd__and3_2 _2980_ (
    .A(\g_bit[6].g_word[24].r_bit.Q ),
    .B(_0297_),
    .C(_0298_),
    .X(_0665_)
  );
  sky130_fd_sc_hd__a2111o_2 _2981_ (
    .A1(\g_bit[6].g_word[29].r_bit.Q ),
    .A2(_0205_),
    .B1(_0663_),
    .C1(_0664_),
    .D1(_0665_),
    .X(_0666_)
  );
  sky130_fd_sc_hd__and3_2 _2982_ (
    .A(\g_bit[6].g_word[27].r_bit.Q ),
    .B(_0220_),
    .C(_0221_),
    .X(_0667_)
  );
  sky130_fd_sc_hd__a221o_2 _2983_ (
    .A1(\g_bit[6].g_word[6].r_bit.Q ),
    .A2(_0216_),
    .B1(_0218_),
    .B2(\g_bit[6].g_word[1].r_bit.Q ),
    .C1(_0667_),
    .X(_0668_)
  );
  sky130_fd_sc_hd__or3_2 _2984_ (
    .A(_0637_),
    .B(_0485_),
    .C(_0230_),
    .X(_0669_)
  );
  sky130_fd_sc_hd__or3_2 _2985_ (
    .A(_0639_),
    .B(_0609_),
    .C(_0232_),
    .X(_0670_)
  );
  sky130_fd_sc_hd__or3_2 _2986_ (
    .A(_0641_),
    .B(_0146_),
    .C(_0141_),
    .X(_0671_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2987_ (
    .A1(_0636_),
    .A2(_0226_),
    .B1(_0669_),
    .C1(_0670_),
    .D1(_0671_),
    .Y(_0672_)
  );
  sky130_fd_sc_hd__buf_1 _2988_ (
    .A(_0174_),
    .X(_0673_)
  );
  sky130_fd_sc_hd__or3_2 _2989_ (
    .A(_0645_),
    .B(_0239_),
    .C(_0673_),
    .X(_0674_)
  );
  sky130_fd_sc_hd__or3_2 _2990_ (
    .A(_0647_),
    .B(_0242_),
    .C(_0166_),
    .X(_0675_)
  );
  sky130_fd_sc_hd__or3_2 _2991_ (
    .A(_0649_),
    .B(_0309_),
    .C(_0148_),
    .X(_0676_)
  );
  sky130_fd_sc_hd__o2111ai_2 _2992_ (
    .A1(_0644_),
    .A2(_0237_),
    .B1(_0674_),
    .C1(_0675_),
    .D1(_0676_),
    .Y(_0677_)
  );
  sky130_fd_sc_hd__or4_2 _2993_ (
    .A(_0666_),
    .B(_0668_),
    .C(_0672_),
    .D(_0677_),
    .X(_0678_)
  );
  sky130_fd_sc_hd__or4_2 _2994_ (
    .A(_0655_),
    .B(_0657_),
    .C(_0662_),
    .D(_0678_),
    .X(_0679_)
  );
  sky130_fd_sc_hd__buf_1 _2995_ (
    .A(_0679_),
    .X(\g_bit[6].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _2996_ (
    .A1(\g_bit[7].g_word[30].r_bit.Q ),
    .A2(_0023_),
    .A3(_0025_),
    .B1(_0030_),
    .B2(\g_bit[7].g_word[28].r_bit.Q ),
    .X(_0680_)
  );
  sky130_fd_sc_hd__a221o_2 _2997_ (
    .A1(\g_bit[7].g_word[4].r_bit.Q ),
    .A2(_0014_),
    .B1(_0021_),
    .B2(\g_bit[7].g_word[26].r_bit.Q ),
    .C1(_0680_),
    .X(_0681_)
  );
  sky130_fd_sc_hd__a22o_2 _2998_ (
    .A1(\g_bit[7].g_word[5].r_bit.Q ),
    .A2(_0043_),
    .B1(_0050_),
    .B2(\g_bit[7].g_word[2].r_bit.Q ),
    .X(_0682_)
  );
  sky130_fd_sc_hd__a221o_2 _2999_ (
    .A1(\g_bit[7].g_word[25].r_bit.Q ),
    .A2(_0035_),
    .B1(_0039_),
    .B2(\g_bit[7].g_word[31].r_bit.Q ),
    .C1(_0682_),
    .X(_0683_)
  );
  sky130_fd_sc_hd__a22o_2 _3000_ (
    .A1(\g_bit[7].g_word[13].r_bit.Q ),
    .A2(_0054_),
    .B1(_0057_),
    .B2(\g_bit[7].g_word[15].r_bit.Q ),
    .X(_0684_)
  );
  sky130_fd_sc_hd__a22o_2 _3001_ (
    .A1(\g_bit[7].g_word[11].r_bit.Q ),
    .A2(_0060_),
    .B1(_0062_),
    .B2(\g_bit[7].g_word[20].r_bit.Q ),
    .X(_0685_)
  );
  sky130_fd_sc_hd__a22o_2 _3002_ (
    .A1(\g_bit[7].g_word[19].r_bit.Q ),
    .A2(_0065_),
    .B1(_0067_),
    .B2(\g_bit[7].g_word[21].r_bit.Q ),
    .X(_0686_)
  );
  sky130_fd_sc_hd__a22o_2 _3003_ (
    .A1(\g_bit[7].g_word[17].r_bit.Q ),
    .A2(_0070_),
    .B1(_0072_),
    .B2(\g_bit[7].g_word[12].r_bit.Q ),
    .X(_0687_)
  );
  sky130_fd_sc_hd__or4_2 _3004_ (
    .A(_0684_),
    .B(_0685_),
    .C(_0686_),
    .D(_0687_),
    .X(_0688_)
  );
  sky130_fd_sc_hd__inv_2 _3005_ (
    .A(\g_bit[7].g_word[7].r_bit.Q ),
    .Y(_0689_)
  );
  sky130_fd_sc_hd__buf_1 _3006_ (
    .A(_0081_),
    .X(_0690_)
  );
  sky130_fd_sc_hd__nor3_2 _3007_ (
    .A(_0689_),
    .B(_0690_),
    .C(_0004_),
    .Y(_0691_)
  );
  sky130_fd_sc_hd__inv_2 _3008_ (
    .A(\g_bit[7].g_word[3].r_bit.Q ),
    .Y(_0692_)
  );
  sky130_fd_sc_hd__nor3_2 _3009_ (
    .A(_0692_),
    .B(_0085_),
    .C(_0086_),
    .Y(_0693_)
  );
  sky130_fd_sc_hd__and3_2 _3010_ (
    .A(\g_bit[7].g_word[24].r_bit.Q ),
    .B(_0260_),
    .C(_0261_),
    .X(_0694_)
  );
  sky130_fd_sc_hd__a2111o_2 _3011_ (
    .A1(\g_bit[7].g_word[29].r_bit.Q ),
    .A2(_0076_),
    .B1(_0691_),
    .C1(_0693_),
    .D1(_0694_),
    .X(_0695_)
  );
  sky130_fd_sc_hd__and3_2 _3012_ (
    .A(\g_bit[7].g_word[27].r_bit.Q ),
    .B(_0094_),
    .C(_0095_),
    .X(_0696_)
  );
  sky130_fd_sc_hd__a221o_2 _3013_ (
    .A1(\g_bit[7].g_word[6].r_bit.Q ),
    .A2(_0090_),
    .B1(_0092_),
    .B2(\g_bit[7].g_word[1].r_bit.Q ),
    .C1(_0696_),
    .X(_0697_)
  );
  sky130_fd_sc_hd__inv_2 _3014_ (
    .A(\g_bit[7].g_word[23].r_bit.Q ),
    .Y(_0698_)
  );
  sky130_fd_sc_hd__inv_2 _3015_ (
    .A(\g_bit[7].g_word[10].r_bit.Q ),
    .Y(_0699_)
  );
  sky130_fd_sc_hd__buf_1 _3016_ (
    .A(_0048_),
    .X(_0700_)
  );
  sky130_fd_sc_hd__or3_2 _3017_ (
    .A(_0699_),
    .B(_0453_),
    .C(_0700_),
    .X(_0701_)
  );
  sky130_fd_sc_hd__inv_2 _3018_ (
    .A(\g_bit[7].g_word[9].r_bit.Q ),
    .Y(_0702_)
  );
  sky130_fd_sc_hd__or3_2 _3019_ (
    .A(_0702_),
    .B(_0577_),
    .C(_0110_),
    .X(_0703_)
  );
  sky130_fd_sc_hd__inv_2 _3020_ (
    .A(\g_bit[7].g_word[8].r_bit.Q ),
    .Y(_0704_)
  );
  sky130_fd_sc_hd__buf_1 _3021_ (
    .A(_0016_),
    .X(_0705_)
  );
  sky130_fd_sc_hd__or3_2 _3022_ (
    .A(_0704_),
    .B(_0705_),
    .C(_0012_),
    .X(_0706_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3023_ (
    .A1(_0698_),
    .A2(_0101_),
    .B1(_0701_),
    .C1(_0703_),
    .D1(_0706_),
    .Y(_0707_)
  );
  sky130_fd_sc_hd__inv_2 _3024_ (
    .A(\g_bit[7].g_word[22].r_bit.Q ),
    .Y(_0708_)
  );
  sky130_fd_sc_hd__inv_2 _3025_ (
    .A(\g_bit[7].g_word[16].r_bit.Q ),
    .Y(_0709_)
  );
  sky130_fd_sc_hd__or3_2 _3026_ (
    .A(_0709_),
    .B(_0584_),
    .C(_0121_),
    .X(_0710_)
  );
  sky130_fd_sc_hd__inv_2 _3027_ (
    .A(\g_bit[7].g_word[14].r_bit.Q ),
    .Y(_0711_)
  );
  sky130_fd_sc_hd__or3_2 _3028_ (
    .A(_0711_),
    .B(_0124_),
    .C(_0037_),
    .X(_0712_)
  );
  sky130_fd_sc_hd__inv_2 _3029_ (
    .A(\g_bit[7].g_word[18].r_bit.Q ),
    .Y(_0713_)
  );
  sky130_fd_sc_hd__or3_2 _3030_ (
    .A(_0713_),
    .B(_0280_),
    .C(_0019_),
    .X(_0714_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3031_ (
    .A1(_0708_),
    .A2(_0116_),
    .B1(_0710_),
    .C1(_0712_),
    .D1(_0714_),
    .Y(_0715_)
  );
  sky130_fd_sc_hd__or4_2 _3032_ (
    .A(_0695_),
    .B(_0697_),
    .C(_0707_),
    .D(_0715_),
    .X(_0716_)
  );
  sky130_fd_sc_hd__or4_2 _3033_ (
    .A(_0681_),
    .B(_0683_),
    .C(_0688_),
    .D(_0716_),
    .X(_0717_)
  );
  sky130_fd_sc_hd__buf_1 _3034_ (
    .A(_0717_),
    .X(\g_bit[7].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _3035_ (
    .A1(\g_bit[7].g_word[30].r_bit.Q ),
    .A2(_0152_),
    .A3(_0154_),
    .B1(_0159_),
    .B2(\g_bit[7].g_word[28].r_bit.Q ),
    .X(_0718_)
  );
  sky130_fd_sc_hd__a221o_2 _3036_ (
    .A1(\g_bit[7].g_word[4].r_bit.Q ),
    .A2(_0143_),
    .B1(_0150_),
    .B2(\g_bit[7].g_word[26].r_bit.Q ),
    .C1(_0718_),
    .X(_0719_)
  );
  sky130_fd_sc_hd__a22o_2 _3037_ (
    .A1(\g_bit[7].g_word[5].r_bit.Q ),
    .A2(_0172_),
    .B1(_0179_),
    .B2(\g_bit[7].g_word[2].r_bit.Q ),
    .X(_0720_)
  );
  sky130_fd_sc_hd__a221o_2 _3038_ (
    .A1(\g_bit[7].g_word[25].r_bit.Q ),
    .A2(_0164_),
    .B1(_0168_),
    .B2(\g_bit[7].g_word[31].r_bit.Q ),
    .C1(_0720_),
    .X(_0721_)
  );
  sky130_fd_sc_hd__a22o_2 _3039_ (
    .A1(\g_bit[7].g_word[13].r_bit.Q ),
    .A2(_0183_),
    .B1(_0186_),
    .B2(\g_bit[7].g_word[15].r_bit.Q ),
    .X(_0722_)
  );
  sky130_fd_sc_hd__a22o_2 _3040_ (
    .A1(\g_bit[7].g_word[20].r_bit.Q ),
    .A2(_0189_),
    .B1(_0191_),
    .B2(\g_bit[7].g_word[11].r_bit.Q ),
    .X(_0723_)
  );
  sky130_fd_sc_hd__a22o_2 _3041_ (
    .A1(\g_bit[7].g_word[19].r_bit.Q ),
    .A2(_0194_),
    .B1(_0196_),
    .B2(\g_bit[7].g_word[21].r_bit.Q ),
    .X(_0724_)
  );
  sky130_fd_sc_hd__a22o_2 _3042_ (
    .A1(\g_bit[7].g_word[17].r_bit.Q ),
    .A2(_0199_),
    .B1(_0201_),
    .B2(\g_bit[7].g_word[12].r_bit.Q ),
    .X(_0725_)
  );
  sky130_fd_sc_hd__or4_2 _3043_ (
    .A(_0722_),
    .B(_0723_),
    .C(_0724_),
    .D(_0725_),
    .X(_0726_)
  );
  sky130_fd_sc_hd__buf_1 _3044_ (
    .A(_0209_),
    .X(_0727_)
  );
  sky130_fd_sc_hd__nor3_2 _3045_ (
    .A(_0689_),
    .B(_0133_),
    .C(_0727_),
    .Y(_0728_)
  );
  sky130_fd_sc_hd__nor3_2 _3046_ (
    .A(_0692_),
    .B(_0212_),
    .C(_0210_),
    .Y(_0729_)
  );
  sky130_fd_sc_hd__and3_2 _3047_ (
    .A(\g_bit[7].g_word[24].r_bit.Q ),
    .B(_0297_),
    .C(_0298_),
    .X(_0730_)
  );
  sky130_fd_sc_hd__a2111o_2 _3048_ (
    .A1(\g_bit[7].g_word[29].r_bit.Q ),
    .A2(_0205_),
    .B1(_0728_),
    .C1(_0729_),
    .D1(_0730_),
    .X(_0731_)
  );
  sky130_fd_sc_hd__and3_2 _3049_ (
    .A(\g_bit[7].g_word[27].r_bit.Q ),
    .B(_0220_),
    .C(_0221_),
    .X(_0732_)
  );
  sky130_fd_sc_hd__a221o_2 _3050_ (
    .A1(\g_bit[7].g_word[6].r_bit.Q ),
    .A2(_0216_),
    .B1(_0218_),
    .B2(\g_bit[7].g_word[1].r_bit.Q ),
    .C1(_0732_),
    .X(_0733_)
  );
  sky130_fd_sc_hd__buf_1 _3051_ (
    .A(_0177_),
    .X(_0734_)
  );
  sky130_fd_sc_hd__or3_2 _3052_ (
    .A(_0699_),
    .B(_0485_),
    .C(_0734_),
    .X(_0735_)
  );
  sky130_fd_sc_hd__or3_2 _3053_ (
    .A(_0702_),
    .B(_0609_),
    .C(_0232_),
    .X(_0736_)
  );
  sky130_fd_sc_hd__buf_1 _3054_ (
    .A(_0145_),
    .X(_0737_)
  );
  sky130_fd_sc_hd__or3_2 _3055_ (
    .A(_0704_),
    .B(_0737_),
    .C(_0141_),
    .X(_0738_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3056_ (
    .A1(_0698_),
    .A2(_0226_),
    .B1(_0735_),
    .C1(_0736_),
    .D1(_0738_),
    .Y(_0739_)
  );
  sky130_fd_sc_hd__or3_2 _3057_ (
    .A(_0709_),
    .B(_0239_),
    .C(_0673_),
    .X(_0740_)
  );
  sky130_fd_sc_hd__or3_2 _3058_ (
    .A(_0711_),
    .B(_0242_),
    .C(_0166_),
    .X(_0741_)
  );
  sky130_fd_sc_hd__or3_2 _3059_ (
    .A(_0713_),
    .B(_0309_),
    .C(_0148_),
    .X(_0742_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3060_ (
    .A1(_0708_),
    .A2(_0237_),
    .B1(_0740_),
    .C1(_0741_),
    .D1(_0742_),
    .Y(_0743_)
  );
  sky130_fd_sc_hd__or4_2 _3061_ (
    .A(_0731_),
    .B(_0733_),
    .C(_0739_),
    .D(_0743_),
    .X(_0744_)
  );
  sky130_fd_sc_hd__or4_2 _3062_ (
    .A(_0719_),
    .B(_0721_),
    .C(_0726_),
    .D(_0744_),
    .X(_0745_)
  );
  sky130_fd_sc_hd__buf_1 _3063_ (
    .A(_0745_),
    .X(\g_bit[7].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _3064_ (
    .A1(\g_bit[8].g_word[30].r_bit.Q ),
    .A2(_0023_),
    .A3(_0025_),
    .B1(_0030_),
    .B2(\g_bit[8].g_word[28].r_bit.Q ),
    .X(_0746_)
  );
  sky130_fd_sc_hd__a221o_2 _3065_ (
    .A1(\g_bit[8].g_word[4].r_bit.Q ),
    .A2(_0014_),
    .B1(_0021_),
    .B2(\g_bit[8].g_word[26].r_bit.Q ),
    .C1(_0746_),
    .X(_0747_)
  );
  sky130_fd_sc_hd__a22o_2 _3066_ (
    .A1(\g_bit[8].g_word[5].r_bit.Q ),
    .A2(_0043_),
    .B1(_0050_),
    .B2(\g_bit[8].g_word[2].r_bit.Q ),
    .X(_0748_)
  );
  sky130_fd_sc_hd__a221o_2 _3067_ (
    .A1(\g_bit[8].g_word[25].r_bit.Q ),
    .A2(_0035_),
    .B1(_0039_),
    .B2(\g_bit[8].g_word[31].r_bit.Q ),
    .C1(_0748_),
    .X(_0749_)
  );
  sky130_fd_sc_hd__a22o_2 _3068_ (
    .A1(\g_bit[8].g_word[13].r_bit.Q ),
    .A2(_0054_),
    .B1(_0057_),
    .B2(\g_bit[8].g_word[15].r_bit.Q ),
    .X(_0750_)
  );
  sky130_fd_sc_hd__a22o_2 _3069_ (
    .A1(\g_bit[8].g_word[11].r_bit.Q ),
    .A2(_0060_),
    .B1(_0062_),
    .B2(\g_bit[8].g_word[20].r_bit.Q ),
    .X(_0751_)
  );
  sky130_fd_sc_hd__a22o_2 _3070_ (
    .A1(\g_bit[8].g_word[19].r_bit.Q ),
    .A2(_0065_),
    .B1(_0067_),
    .B2(\g_bit[8].g_word[21].r_bit.Q ),
    .X(_0752_)
  );
  sky130_fd_sc_hd__a22o_2 _3071_ (
    .A1(\g_bit[8].g_word[17].r_bit.Q ),
    .A2(_0070_),
    .B1(_0072_),
    .B2(\g_bit[8].g_word[12].r_bit.Q ),
    .X(_0753_)
  );
  sky130_fd_sc_hd__or4_2 _3072_ (
    .A(_0750_),
    .B(_0751_),
    .C(_0752_),
    .D(_0753_),
    .X(_0754_)
  );
  sky130_fd_sc_hd__inv_2 _3073_ (
    .A(\g_bit[8].g_word[7].r_bit.Q ),
    .Y(_0755_)
  );
  sky130_fd_sc_hd__buf_1 _3074_ (
    .A(_0003_),
    .X(_0756_)
  );
  sky130_fd_sc_hd__nor3_2 _3075_ (
    .A(_0755_),
    .B(_0690_),
    .C(_0756_),
    .Y(_0757_)
  );
  sky130_fd_sc_hd__inv_2 _3076_ (
    .A(\g_bit[8].g_word[3].r_bit.Q ),
    .Y(_0758_)
  );
  sky130_fd_sc_hd__nor3_2 _3077_ (
    .A(_0758_),
    .B(_0085_),
    .C(_0086_),
    .Y(_0759_)
  );
  sky130_fd_sc_hd__buf_1 _3078_ (
    .A(_0077_),
    .X(_0760_)
  );
  sky130_fd_sc_hd__and3_2 _3079_ (
    .A(\g_bit[8].g_word[24].r_bit.Q ),
    .B(_0760_),
    .C(_0261_),
    .X(_0761_)
  );
  sky130_fd_sc_hd__a2111o_2 _3080_ (
    .A1(\g_bit[8].g_word[29].r_bit.Q ),
    .A2(_0076_),
    .B1(_0757_),
    .C1(_0759_),
    .D1(_0761_),
    .X(_0762_)
  );
  sky130_fd_sc_hd__and3_2 _3081_ (
    .A(\g_bit[8].g_word[27].r_bit.Q ),
    .B(_0094_),
    .C(_0095_),
    .X(_0763_)
  );
  sky130_fd_sc_hd__a221o_2 _3082_ (
    .A1(\g_bit[8].g_word[6].r_bit.Q ),
    .A2(_0090_),
    .B1(_0092_),
    .B2(\g_bit[8].g_word[1].r_bit.Q ),
    .C1(_0763_),
    .X(_0764_)
  );
  sky130_fd_sc_hd__inv_2 _3083_ (
    .A(\g_bit[8].g_word[23].r_bit.Q ),
    .Y(_0765_)
  );
  sky130_fd_sc_hd__inv_2 _3084_ (
    .A(\g_bit[8].g_word[10].r_bit.Q ),
    .Y(_0766_)
  );
  sky130_fd_sc_hd__or3_2 _3085_ (
    .A(_0766_),
    .B(_0453_),
    .C(_0700_),
    .X(_0767_)
  );
  sky130_fd_sc_hd__inv_2 _3086_ (
    .A(\g_bit[8].g_word[9].r_bit.Q ),
    .Y(_0768_)
  );
  sky130_fd_sc_hd__or3_2 _3087_ (
    .A(_0768_),
    .B(_0577_),
    .C(_0110_),
    .X(_0769_)
  );
  sky130_fd_sc_hd__inv_2 _3088_ (
    .A(\g_bit[8].g_word[8].r_bit.Q ),
    .Y(_0770_)
  );
  sky130_fd_sc_hd__or3_2 _3089_ (
    .A(_0770_),
    .B(_0705_),
    .C(_0012_),
    .X(_0771_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3090_ (
    .A1(_0765_),
    .A2(_0101_),
    .B1(_0767_),
    .C1(_0769_),
    .D1(_0771_),
    .Y(_0772_)
  );
  sky130_fd_sc_hd__inv_2 _3091_ (
    .A(\g_bit[8].g_word[22].r_bit.Q ),
    .Y(_0773_)
  );
  sky130_fd_sc_hd__inv_2 _3092_ (
    .A(\g_bit[8].g_word[16].r_bit.Q ),
    .Y(_0774_)
  );
  sky130_fd_sc_hd__or3_2 _3093_ (
    .A(_0774_),
    .B(_0584_),
    .C(_0121_),
    .X(_0775_)
  );
  sky130_fd_sc_hd__inv_2 _3094_ (
    .A(\g_bit[8].g_word[14].r_bit.Q ),
    .Y(_0776_)
  );
  sky130_fd_sc_hd__buf_1 _3095_ (
    .A(_0028_),
    .X(_0777_)
  );
  sky130_fd_sc_hd__or3_2 _3096_ (
    .A(_0776_),
    .B(_0124_),
    .C(_0777_),
    .X(_0778_)
  );
  sky130_fd_sc_hd__inv_2 _3097_ (
    .A(\g_bit[8].g_word[18].r_bit.Q ),
    .Y(_0779_)
  );
  sky130_fd_sc_hd__buf_1 _3098_ (
    .A(_0046_),
    .X(_0780_)
  );
  sky130_fd_sc_hd__or3_2 _3099_ (
    .A(_0779_),
    .B(_0780_),
    .C(_0019_),
    .X(_0781_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3100_ (
    .A1(_0773_),
    .A2(_0116_),
    .B1(_0775_),
    .C1(_0778_),
    .D1(_0781_),
    .Y(_0782_)
  );
  sky130_fd_sc_hd__or4_2 _3101_ (
    .A(_0762_),
    .B(_0764_),
    .C(_0772_),
    .D(_0782_),
    .X(_0783_)
  );
  sky130_fd_sc_hd__or4_2 _3102_ (
    .A(_0747_),
    .B(_0749_),
    .C(_0754_),
    .D(_0783_),
    .X(_0784_)
  );
  sky130_fd_sc_hd__buf_1 _3103_ (
    .A(_0784_),
    .X(\g_bit[8].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _3104_ (
    .A1(\g_bit[8].g_word[30].r_bit.Q ),
    .A2(_0152_),
    .A3(_0154_),
    .B1(_0159_),
    .B2(\g_bit[8].g_word[28].r_bit.Q ),
    .X(_0785_)
  );
  sky130_fd_sc_hd__a221o_2 _3105_ (
    .A1(\g_bit[8].g_word[4].r_bit.Q ),
    .A2(_0143_),
    .B1(_0150_),
    .B2(\g_bit[8].g_word[26].r_bit.Q ),
    .C1(_0785_),
    .X(_0786_)
  );
  sky130_fd_sc_hd__a22o_2 _3106_ (
    .A1(\g_bit[8].g_word[5].r_bit.Q ),
    .A2(_0172_),
    .B1(_0179_),
    .B2(\g_bit[8].g_word[2].r_bit.Q ),
    .X(_0787_)
  );
  sky130_fd_sc_hd__a221o_2 _3107_ (
    .A1(\g_bit[8].g_word[25].r_bit.Q ),
    .A2(_0164_),
    .B1(_0168_),
    .B2(\g_bit[8].g_word[31].r_bit.Q ),
    .C1(_0787_),
    .X(_0788_)
  );
  sky130_fd_sc_hd__a22o_2 _3108_ (
    .A1(\g_bit[8].g_word[13].r_bit.Q ),
    .A2(_0183_),
    .B1(_0186_),
    .B2(\g_bit[8].g_word[15].r_bit.Q ),
    .X(_0789_)
  );
  sky130_fd_sc_hd__a22o_2 _3109_ (
    .A1(\g_bit[8].g_word[20].r_bit.Q ),
    .A2(_0189_),
    .B1(_0191_),
    .B2(\g_bit[8].g_word[11].r_bit.Q ),
    .X(_0790_)
  );
  sky130_fd_sc_hd__a22o_2 _3110_ (
    .A1(\g_bit[8].g_word[19].r_bit.Q ),
    .A2(_0194_),
    .B1(_0196_),
    .B2(\g_bit[8].g_word[21].r_bit.Q ),
    .X(_0791_)
  );
  sky130_fd_sc_hd__a22o_2 _3111_ (
    .A1(\g_bit[8].g_word[17].r_bit.Q ),
    .A2(_0199_),
    .B1(_0201_),
    .B2(\g_bit[8].g_word[12].r_bit.Q ),
    .X(_0792_)
  );
  sky130_fd_sc_hd__or4_2 _3112_ (
    .A(_0789_),
    .B(_0790_),
    .C(_0791_),
    .D(_0792_),
    .X(_0793_)
  );
  sky130_fd_sc_hd__buf_1 _3113_ (
    .A(_0132_),
    .X(_0794_)
  );
  sky130_fd_sc_hd__nor3_2 _3114_ (
    .A(_0755_),
    .B(_0794_),
    .C(_0727_),
    .Y(_0795_)
  );
  sky130_fd_sc_hd__buf_1 _3115_ (
    .A(_0209_),
    .X(_0796_)
  );
  sky130_fd_sc_hd__nor3_2 _3116_ (
    .A(_0758_),
    .B(_0212_),
    .C(_0796_),
    .Y(_0797_)
  );
  sky130_fd_sc_hd__buf_1 _3117_ (
    .A(_0207_),
    .X(_0798_)
  );
  sky130_fd_sc_hd__and3_2 _3118_ (
    .A(\g_bit[8].g_word[24].r_bit.Q ),
    .B(_0297_),
    .C(_0798_),
    .X(_0799_)
  );
  sky130_fd_sc_hd__a2111o_2 _3119_ (
    .A1(\g_bit[8].g_word[29].r_bit.Q ),
    .A2(_0205_),
    .B1(_0795_),
    .C1(_0797_),
    .D1(_0799_),
    .X(_0800_)
  );
  sky130_fd_sc_hd__and3_2 _3120_ (
    .A(\g_bit[8].g_word[27].r_bit.Q ),
    .B(_0220_),
    .C(_0221_),
    .X(_0801_)
  );
  sky130_fd_sc_hd__a221o_2 _3121_ (
    .A1(\g_bit[8].g_word[6].r_bit.Q ),
    .A2(_0216_),
    .B1(_0218_),
    .B2(\g_bit[8].g_word[1].r_bit.Q ),
    .C1(_0801_),
    .X(_0802_)
  );
  sky130_fd_sc_hd__or3_2 _3122_ (
    .A(_0766_),
    .B(_0485_),
    .C(_0734_),
    .X(_0803_)
  );
  sky130_fd_sc_hd__or3_2 _3123_ (
    .A(_0768_),
    .B(_0609_),
    .C(_0232_),
    .X(_0804_)
  );
  sky130_fd_sc_hd__or3_2 _3124_ (
    .A(_0770_),
    .B(_0737_),
    .C(_0141_),
    .X(_0805_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3125_ (
    .A1(_0765_),
    .A2(_0226_),
    .B1(_0803_),
    .C1(_0804_),
    .D1(_0805_),
    .Y(_0806_)
  );
  sky130_fd_sc_hd__or3_2 _3126_ (
    .A(_0774_),
    .B(_0239_),
    .C(_0673_),
    .X(_0807_)
  );
  sky130_fd_sc_hd__buf_1 _3127_ (
    .A(_0157_),
    .X(_0808_)
  );
  sky130_fd_sc_hd__or3_2 _3128_ (
    .A(_0776_),
    .B(_0242_),
    .C(_0808_),
    .X(_0809_)
  );
  sky130_fd_sc_hd__buf_1 _3129_ (
    .A(_0175_),
    .X(_0810_)
  );
  sky130_fd_sc_hd__or3_2 _3130_ (
    .A(_0779_),
    .B(_0810_),
    .C(_0148_),
    .X(_0811_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3131_ (
    .A1(_0773_),
    .A2(_0237_),
    .B1(_0807_),
    .C1(_0809_),
    .D1(_0811_),
    .Y(_0812_)
  );
  sky130_fd_sc_hd__or4_2 _3132_ (
    .A(_0800_),
    .B(_0802_),
    .C(_0806_),
    .D(_0812_),
    .X(_0813_)
  );
  sky130_fd_sc_hd__or4_2 _3133_ (
    .A(_0786_),
    .B(_0788_),
    .C(_0793_),
    .D(_0813_),
    .X(_0814_)
  );
  sky130_fd_sc_hd__buf_1 _3134_ (
    .A(_0814_),
    .X(\g_bit[8].r_rs2.D )
  );
  sky130_fd_sc_hd__buf_1 _3135_ (
    .A(_0013_),
    .X(_0815_)
  );
  sky130_fd_sc_hd__buf_1 _3136_ (
    .A(_0020_),
    .X(_0816_)
  );
  sky130_fd_sc_hd__buf_1 _3137_ (
    .A(_0022_),
    .X(_0817_)
  );
  sky130_fd_sc_hd__buf_1 _3138_ (
    .A(_0024_),
    .X(_0818_)
  );
  sky130_fd_sc_hd__buf_1 _3139_ (
    .A(_0029_),
    .X(_0819_)
  );
  sky130_fd_sc_hd__a32o_2 _3140_ (
    .A1(\g_bit[9].g_word[30].r_bit.Q ),
    .A2(_0817_),
    .A3(_0818_),
    .B1(_0819_),
    .B2(\g_bit[9].g_word[28].r_bit.Q ),
    .X(_0820_)
  );
  sky130_fd_sc_hd__a221o_2 _3141_ (
    .A1(\g_bit[9].g_word[4].r_bit.Q ),
    .A2(_0815_),
    .B1(_0816_),
    .B2(\g_bit[9].g_word[26].r_bit.Q ),
    .C1(_0820_),
    .X(_0821_)
  );
  sky130_fd_sc_hd__buf_1 _3142_ (
    .A(_0034_),
    .X(_0822_)
  );
  sky130_fd_sc_hd__buf_1 _3143_ (
    .A(_0038_),
    .X(_0823_)
  );
  sky130_fd_sc_hd__buf_1 _3144_ (
    .A(_0042_),
    .X(_0824_)
  );
  sky130_fd_sc_hd__buf_1 _3145_ (
    .A(_0049_),
    .X(_0825_)
  );
  sky130_fd_sc_hd__a22o_2 _3146_ (
    .A1(\g_bit[9].g_word[5].r_bit.Q ),
    .A2(_0824_),
    .B1(_0825_),
    .B2(\g_bit[9].g_word[2].r_bit.Q ),
    .X(_0826_)
  );
  sky130_fd_sc_hd__a221o_2 _3147_ (
    .A1(\g_bit[9].g_word[25].r_bit.Q ),
    .A2(_0822_),
    .B1(_0823_),
    .B2(\g_bit[9].g_word[31].r_bit.Q ),
    .C1(_0826_),
    .X(_0827_)
  );
  sky130_fd_sc_hd__buf_1 _3148_ (
    .A(_0053_),
    .X(_0828_)
  );
  sky130_fd_sc_hd__buf_1 _3149_ (
    .A(_0056_),
    .X(_0829_)
  );
  sky130_fd_sc_hd__a22o_2 _3150_ (
    .A1(\g_bit[9].g_word[13].r_bit.Q ),
    .A2(_0828_),
    .B1(_0829_),
    .B2(\g_bit[9].g_word[15].r_bit.Q ),
    .X(_0830_)
  );
  sky130_fd_sc_hd__buf_1 _3151_ (
    .A(_0059_),
    .X(_0831_)
  );
  sky130_fd_sc_hd__buf_1 _3152_ (
    .A(_0061_),
    .X(_0832_)
  );
  sky130_fd_sc_hd__a22o_2 _3153_ (
    .A1(\g_bit[9].g_word[11].r_bit.Q ),
    .A2(_0831_),
    .B1(_0832_),
    .B2(\g_bit[9].g_word[20].r_bit.Q ),
    .X(_0833_)
  );
  sky130_fd_sc_hd__buf_1 _3154_ (
    .A(_0064_),
    .X(_0834_)
  );
  sky130_fd_sc_hd__buf_1 _3155_ (
    .A(_0066_),
    .X(_0835_)
  );
  sky130_fd_sc_hd__a22o_2 _3156_ (
    .A1(\g_bit[9].g_word[19].r_bit.Q ),
    .A2(_0834_),
    .B1(_0835_),
    .B2(\g_bit[9].g_word[21].r_bit.Q ),
    .X(_0836_)
  );
  sky130_fd_sc_hd__buf_1 _3157_ (
    .A(_0069_),
    .X(_0837_)
  );
  sky130_fd_sc_hd__buf_1 _3158_ (
    .A(_0071_),
    .X(_0838_)
  );
  sky130_fd_sc_hd__a22o_2 _3159_ (
    .A1(\g_bit[9].g_word[17].r_bit.Q ),
    .A2(_0837_),
    .B1(_0838_),
    .B2(\g_bit[9].g_word[12].r_bit.Q ),
    .X(_0839_)
  );
  sky130_fd_sc_hd__or4_2 _3160_ (
    .A(_0830_),
    .B(_0833_),
    .C(_0836_),
    .D(_0839_),
    .X(_0840_)
  );
  sky130_fd_sc_hd__buf_1 _3161_ (
    .A(_0075_),
    .X(_0841_)
  );
  sky130_fd_sc_hd__inv_2 _3162_ (
    .A(\g_bit[9].g_word[7].r_bit.Q ),
    .Y(_0842_)
  );
  sky130_fd_sc_hd__nor3_2 _3163_ (
    .A(_0842_),
    .B(_0690_),
    .C(_0756_),
    .Y(_0843_)
  );
  sky130_fd_sc_hd__inv_2 _3164_ (
    .A(\g_bit[9].g_word[3].r_bit.Q ),
    .Y(_0844_)
  );
  sky130_fd_sc_hd__buf_1 _3165_ (
    .A(_0045_),
    .X(_0845_)
  );
  sky130_fd_sc_hd__buf_1 _3166_ (
    .A(_0081_),
    .X(_0846_)
  );
  sky130_fd_sc_hd__nor3_2 _3167_ (
    .A(_0844_),
    .B(_0845_),
    .C(_0846_),
    .Y(_0847_)
  );
  sky130_fd_sc_hd__and3_2 _3168_ (
    .A(\g_bit[9].g_word[24].r_bit.Q ),
    .B(_0760_),
    .C(_0261_),
    .X(_0848_)
  );
  sky130_fd_sc_hd__a2111o_2 _3169_ (
    .A1(\g_bit[9].g_word[29].r_bit.Q ),
    .A2(_0841_),
    .B1(_0843_),
    .C1(_0847_),
    .D1(_0848_),
    .X(_0849_)
  );
  sky130_fd_sc_hd__buf_1 _3170_ (
    .A(_0089_),
    .X(_0850_)
  );
  sky130_fd_sc_hd__buf_1 _3171_ (
    .A(_0091_),
    .X(_0851_)
  );
  sky130_fd_sc_hd__buf_1 _3172_ (
    .A(_0093_),
    .X(_0852_)
  );
  sky130_fd_sc_hd__buf_1 _3173_ (
    .A(_0077_),
    .X(_0853_)
  );
  sky130_fd_sc_hd__and3_2 _3174_ (
    .A(\g_bit[9].g_word[27].r_bit.Q ),
    .B(_0852_),
    .C(_0853_),
    .X(_0854_)
  );
  sky130_fd_sc_hd__a221o_2 _3175_ (
    .A1(\g_bit[9].g_word[6].r_bit.Q ),
    .A2(_0850_),
    .B1(_0851_),
    .B2(\g_bit[9].g_word[1].r_bit.Q ),
    .C1(_0854_),
    .X(_0855_)
  );
  sky130_fd_sc_hd__inv_2 _3176_ (
    .A(\g_bit[9].g_word[23].r_bit.Q ),
    .Y(_0856_)
  );
  sky130_fd_sc_hd__buf_1 _3177_ (
    .A(_0100_),
    .X(_0857_)
  );
  sky130_fd_sc_hd__inv_2 _3178_ (
    .A(\g_bit[9].g_word[10].r_bit.Q ),
    .Y(_0858_)
  );
  sky130_fd_sc_hd__or3_2 _3179_ (
    .A(_0858_),
    .B(_0453_),
    .C(_0700_),
    .X(_0859_)
  );
  sky130_fd_sc_hd__inv_2 _3180_ (
    .A(\g_bit[9].g_word[9].r_bit.Q ),
    .Y(_0860_)
  );
  sky130_fd_sc_hd__buf_1 _3181_ (
    .A(_0041_),
    .X(_0861_)
  );
  sky130_fd_sc_hd__or3_2 _3182_ (
    .A(_0860_),
    .B(_0577_),
    .C(_0861_),
    .X(_0862_)
  );
  sky130_fd_sc_hd__inv_2 _3183_ (
    .A(\g_bit[9].g_word[8].r_bit.Q ),
    .Y(_0863_)
  );
  sky130_fd_sc_hd__buf_1 _3184_ (
    .A(_0011_),
    .X(_0864_)
  );
  sky130_fd_sc_hd__or3_2 _3185_ (
    .A(_0863_),
    .B(_0705_),
    .C(_0864_),
    .X(_0865_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3186_ (
    .A1(_0856_),
    .A2(_0857_),
    .B1(_0859_),
    .C1(_0862_),
    .D1(_0865_),
    .Y(_0866_)
  );
  sky130_fd_sc_hd__inv_2 _3187_ (
    .A(\g_bit[9].g_word[22].r_bit.Q ),
    .Y(_0867_)
  );
  sky130_fd_sc_hd__buf_1 _3188_ (
    .A(_0115_),
    .X(_0868_)
  );
  sky130_fd_sc_hd__inv_2 _3189_ (
    .A(\g_bit[9].g_word[16].r_bit.Q ),
    .Y(_0869_)
  );
  sky130_fd_sc_hd__buf_1 _3190_ (
    .A(_0026_),
    .X(_0870_)
  );
  sky130_fd_sc_hd__or3_2 _3191_ (
    .A(_0869_),
    .B(_0584_),
    .C(_0870_),
    .X(_0871_)
  );
  sky130_fd_sc_hd__inv_2 _3192_ (
    .A(\g_bit[9].g_word[14].r_bit.Q ),
    .Y(_0872_)
  );
  sky130_fd_sc_hd__buf_1 _3193_ (
    .A(_0048_),
    .X(_0873_)
  );
  sky130_fd_sc_hd__or3_2 _3194_ (
    .A(_0872_),
    .B(_0873_),
    .C(_0777_),
    .X(_0874_)
  );
  sky130_fd_sc_hd__inv_2 _3195_ (
    .A(\g_bit[9].g_word[18].r_bit.Q ),
    .Y(_0875_)
  );
  sky130_fd_sc_hd__buf_1 _3196_ (
    .A(_0018_),
    .X(_0876_)
  );
  sky130_fd_sc_hd__or3_2 _3197_ (
    .A(_0875_),
    .B(_0780_),
    .C(_0876_),
    .X(_0877_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3198_ (
    .A1(_0867_),
    .A2(_0868_),
    .B1(_0871_),
    .C1(_0874_),
    .D1(_0877_),
    .Y(_0878_)
  );
  sky130_fd_sc_hd__or4_2 _3199_ (
    .A(_0849_),
    .B(_0855_),
    .C(_0866_),
    .D(_0878_),
    .X(_0879_)
  );
  sky130_fd_sc_hd__or4_2 _3200_ (
    .A(_0821_),
    .B(_0827_),
    .C(_0840_),
    .D(_0879_),
    .X(_0880_)
  );
  sky130_fd_sc_hd__buf_1 _3201_ (
    .A(_0880_),
    .X(\g_bit[9].r_rs1.D )
  );
  sky130_fd_sc_hd__buf_1 _3202_ (
    .A(_0142_),
    .X(_0881_)
  );
  sky130_fd_sc_hd__buf_1 _3203_ (
    .A(_0149_),
    .X(_0882_)
  );
  sky130_fd_sc_hd__buf_1 _3204_ (
    .A(_0151_),
    .X(_0883_)
  );
  sky130_fd_sc_hd__buf_1 _3205_ (
    .A(_0153_),
    .X(_0884_)
  );
  sky130_fd_sc_hd__buf_1 _3206_ (
    .A(_0158_),
    .X(_0885_)
  );
  sky130_fd_sc_hd__a32o_2 _3207_ (
    .A1(\g_bit[9].g_word[30].r_bit.Q ),
    .A2(_0883_),
    .A3(_0884_),
    .B1(_0885_),
    .B2(\g_bit[9].g_word[28].r_bit.Q ),
    .X(_0886_)
  );
  sky130_fd_sc_hd__a221o_2 _3208_ (
    .A1(\g_bit[9].g_word[4].r_bit.Q ),
    .A2(_0881_),
    .B1(_0882_),
    .B2(\g_bit[9].g_word[26].r_bit.Q ),
    .C1(_0886_),
    .X(_0887_)
  );
  sky130_fd_sc_hd__buf_1 _3209_ (
    .A(_0163_),
    .X(_0888_)
  );
  sky130_fd_sc_hd__buf_1 _3210_ (
    .A(_0167_),
    .X(_0889_)
  );
  sky130_fd_sc_hd__buf_1 _3211_ (
    .A(_0171_),
    .X(_0890_)
  );
  sky130_fd_sc_hd__buf_1 _3212_ (
    .A(_0178_),
    .X(_0891_)
  );
  sky130_fd_sc_hd__a22o_2 _3213_ (
    .A1(\g_bit[9].g_word[5].r_bit.Q ),
    .A2(_0890_),
    .B1(_0891_),
    .B2(\g_bit[9].g_word[2].r_bit.Q ),
    .X(_0892_)
  );
  sky130_fd_sc_hd__a221o_2 _3214_ (
    .A1(\g_bit[9].g_word[25].r_bit.Q ),
    .A2(_0888_),
    .B1(_0889_),
    .B2(\g_bit[9].g_word[31].r_bit.Q ),
    .C1(_0892_),
    .X(_0893_)
  );
  sky130_fd_sc_hd__buf_1 _3215_ (
    .A(_0182_),
    .X(_0894_)
  );
  sky130_fd_sc_hd__buf_1 _3216_ (
    .A(_0185_),
    .X(_0895_)
  );
  sky130_fd_sc_hd__a22o_2 _3217_ (
    .A1(\g_bit[9].g_word[13].r_bit.Q ),
    .A2(_0894_),
    .B1(_0895_),
    .B2(\g_bit[9].g_word[15].r_bit.Q ),
    .X(_0896_)
  );
  sky130_fd_sc_hd__buf_1 _3218_ (
    .A(_0188_),
    .X(_0897_)
  );
  sky130_fd_sc_hd__buf_1 _3219_ (
    .A(_0190_),
    .X(_0898_)
  );
  sky130_fd_sc_hd__a22o_2 _3220_ (
    .A1(\g_bit[9].g_word[20].r_bit.Q ),
    .A2(_0897_),
    .B1(_0898_),
    .B2(\g_bit[9].g_word[11].r_bit.Q ),
    .X(_0899_)
  );
  sky130_fd_sc_hd__buf_1 _3221_ (
    .A(_0193_),
    .X(_0900_)
  );
  sky130_fd_sc_hd__buf_1 _3222_ (
    .A(_0195_),
    .X(_0901_)
  );
  sky130_fd_sc_hd__a22o_2 _3223_ (
    .A1(\g_bit[9].g_word[19].r_bit.Q ),
    .A2(_0900_),
    .B1(_0901_),
    .B2(\g_bit[9].g_word[21].r_bit.Q ),
    .X(_0902_)
  );
  sky130_fd_sc_hd__buf_1 _3224_ (
    .A(_0198_),
    .X(_0903_)
  );
  sky130_fd_sc_hd__buf_1 _3225_ (
    .A(_0200_),
    .X(_0904_)
  );
  sky130_fd_sc_hd__a22o_2 _3226_ (
    .A1(\g_bit[9].g_word[17].r_bit.Q ),
    .A2(_0903_),
    .B1(_0904_),
    .B2(\g_bit[9].g_word[12].r_bit.Q ),
    .X(_0905_)
  );
  sky130_fd_sc_hd__or4_2 _3227_ (
    .A(_0896_),
    .B(_0899_),
    .C(_0902_),
    .D(_0905_),
    .X(_0906_)
  );
  sky130_fd_sc_hd__buf_1 _3228_ (
    .A(_0204_),
    .X(_0907_)
  );
  sky130_fd_sc_hd__nor3_2 _3229_ (
    .A(_0842_),
    .B(_0794_),
    .C(_0727_),
    .Y(_0908_)
  );
  sky130_fd_sc_hd__buf_1 _3230_ (
    .A(_0174_),
    .X(_0909_)
  );
  sky130_fd_sc_hd__nor3_2 _3231_ (
    .A(_0844_),
    .B(_0909_),
    .C(_0796_),
    .Y(_0910_)
  );
  sky130_fd_sc_hd__and3_2 _3232_ (
    .A(\g_bit[9].g_word[24].r_bit.Q ),
    .B(_0297_),
    .C(_0798_),
    .X(_0911_)
  );
  sky130_fd_sc_hd__a2111o_2 _3233_ (
    .A1(\g_bit[9].g_word[29].r_bit.Q ),
    .A2(_0907_),
    .B1(_0908_),
    .C1(_0910_),
    .D1(_0911_),
    .X(_0912_)
  );
  sky130_fd_sc_hd__buf_1 _3234_ (
    .A(_0215_),
    .X(_0913_)
  );
  sky130_fd_sc_hd__buf_1 _3235_ (
    .A(_0217_),
    .X(_0914_)
  );
  sky130_fd_sc_hd__buf_1 _3236_ (
    .A(_0219_),
    .X(_0915_)
  );
  sky130_fd_sc_hd__buf_1 _3237_ (
    .A(_0207_),
    .X(_0916_)
  );
  sky130_fd_sc_hd__and3_2 _3238_ (
    .A(\g_bit[9].g_word[27].r_bit.Q ),
    .B(_0915_),
    .C(_0916_),
    .X(_0917_)
  );
  sky130_fd_sc_hd__a221o_2 _3239_ (
    .A1(\g_bit[9].g_word[6].r_bit.Q ),
    .A2(_0913_),
    .B1(_0914_),
    .B2(\g_bit[9].g_word[1].r_bit.Q ),
    .C1(_0917_),
    .X(_0918_)
  );
  sky130_fd_sc_hd__buf_1 _3240_ (
    .A(_0225_),
    .X(_0919_)
  );
  sky130_fd_sc_hd__or3_2 _3241_ (
    .A(_0858_),
    .B(_0485_),
    .C(_0734_),
    .X(_0920_)
  );
  sky130_fd_sc_hd__buf_1 _3242_ (
    .A(_0170_),
    .X(_0921_)
  );
  sky130_fd_sc_hd__or3_2 _3243_ (
    .A(_0860_),
    .B(_0609_),
    .C(_0921_),
    .X(_0922_)
  );
  sky130_fd_sc_hd__buf_1 _3244_ (
    .A(_0140_),
    .X(_0923_)
  );
  sky130_fd_sc_hd__or3_2 _3245_ (
    .A(_0863_),
    .B(_0737_),
    .C(_0923_),
    .X(_0924_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3246_ (
    .A1(_0856_),
    .A2(_0919_),
    .B1(_0920_),
    .C1(_0922_),
    .D1(_0924_),
    .Y(_0925_)
  );
  sky130_fd_sc_hd__buf_1 _3247_ (
    .A(_0236_),
    .X(_0926_)
  );
  sky130_fd_sc_hd__buf_1 _3248_ (
    .A(_0155_),
    .X(_0927_)
  );
  sky130_fd_sc_hd__or3_2 _3249_ (
    .A(_0869_),
    .B(_0927_),
    .C(_0673_),
    .X(_0928_)
  );
  sky130_fd_sc_hd__buf_1 _3250_ (
    .A(_0177_),
    .X(_0929_)
  );
  sky130_fd_sc_hd__or3_2 _3251_ (
    .A(_0872_),
    .B(_0929_),
    .C(_0808_),
    .X(_0930_)
  );
  sky130_fd_sc_hd__buf_1 _3252_ (
    .A(_0147_),
    .X(_0931_)
  );
  sky130_fd_sc_hd__or3_2 _3253_ (
    .A(_0875_),
    .B(_0810_),
    .C(_0931_),
    .X(_0932_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3254_ (
    .A1(_0867_),
    .A2(_0926_),
    .B1(_0928_),
    .C1(_0930_),
    .D1(_0932_),
    .Y(_0933_)
  );
  sky130_fd_sc_hd__or4_2 _3255_ (
    .A(_0912_),
    .B(_0918_),
    .C(_0925_),
    .D(_0933_),
    .X(_0934_)
  );
  sky130_fd_sc_hd__or4_2 _3256_ (
    .A(_0887_),
    .B(_0893_),
    .C(_0906_),
    .D(_0934_),
    .X(_0935_)
  );
  sky130_fd_sc_hd__buf_1 _3257_ (
    .A(_0935_),
    .X(\g_bit[9].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _3258_ (
    .A1(\g_bit[10].g_word[30].r_bit.Q ),
    .A2(_0817_),
    .A3(_0818_),
    .B1(_0819_),
    .B2(\g_bit[10].g_word[28].r_bit.Q ),
    .X(_0936_)
  );
  sky130_fd_sc_hd__a221o_2 _3259_ (
    .A1(\g_bit[10].g_word[4].r_bit.Q ),
    .A2(_0815_),
    .B1(_0816_),
    .B2(\g_bit[10].g_word[26].r_bit.Q ),
    .C1(_0936_),
    .X(_0937_)
  );
  sky130_fd_sc_hd__a22o_2 _3260_ (
    .A1(\g_bit[10].g_word[5].r_bit.Q ),
    .A2(_0824_),
    .B1(_0825_),
    .B2(\g_bit[10].g_word[2].r_bit.Q ),
    .X(_0938_)
  );
  sky130_fd_sc_hd__a221o_2 _3261_ (
    .A1(\g_bit[10].g_word[25].r_bit.Q ),
    .A2(_0822_),
    .B1(_0823_),
    .B2(\g_bit[10].g_word[31].r_bit.Q ),
    .C1(_0938_),
    .X(_0939_)
  );
  sky130_fd_sc_hd__a22o_2 _3262_ (
    .A1(\g_bit[10].g_word[13].r_bit.Q ),
    .A2(_0828_),
    .B1(_0829_),
    .B2(\g_bit[10].g_word[15].r_bit.Q ),
    .X(_0940_)
  );
  sky130_fd_sc_hd__a22o_2 _3263_ (
    .A1(\g_bit[10].g_word[11].r_bit.Q ),
    .A2(_0831_),
    .B1(_0832_),
    .B2(\g_bit[10].g_word[20].r_bit.Q ),
    .X(_0941_)
  );
  sky130_fd_sc_hd__a22o_2 _3264_ (
    .A1(\g_bit[10].g_word[19].r_bit.Q ),
    .A2(_0834_),
    .B1(_0835_),
    .B2(\g_bit[10].g_word[21].r_bit.Q ),
    .X(_0942_)
  );
  sky130_fd_sc_hd__a22o_2 _3265_ (
    .A1(\g_bit[10].g_word[17].r_bit.Q ),
    .A2(_0837_),
    .B1(_0838_),
    .B2(\g_bit[10].g_word[12].r_bit.Q ),
    .X(_0943_)
  );
  sky130_fd_sc_hd__or4_2 _3266_ (
    .A(_0940_),
    .B(_0941_),
    .C(_0942_),
    .D(_0943_),
    .X(_0944_)
  );
  sky130_fd_sc_hd__inv_2 _3267_ (
    .A(\g_bit[10].g_word[7].r_bit.Q ),
    .Y(_0945_)
  );
  sky130_fd_sc_hd__nor3_2 _3268_ (
    .A(_0945_),
    .B(_0690_),
    .C(_0756_),
    .Y(_0946_)
  );
  sky130_fd_sc_hd__inv_2 _3269_ (
    .A(\g_bit[10].g_word[3].r_bit.Q ),
    .Y(_0947_)
  );
  sky130_fd_sc_hd__nor3_2 _3270_ (
    .A(_0947_),
    .B(_0845_),
    .C(_0846_),
    .Y(_0948_)
  );
  sky130_fd_sc_hd__buf_1 _3271_ (
    .A(_0078_),
    .X(_0949_)
  );
  sky130_fd_sc_hd__and3_2 _3272_ (
    .A(\g_bit[10].g_word[24].r_bit.Q ),
    .B(_0760_),
    .C(_0949_),
    .X(_0950_)
  );
  sky130_fd_sc_hd__a2111o_2 _3273_ (
    .A1(\g_bit[10].g_word[29].r_bit.Q ),
    .A2(_0841_),
    .B1(_0946_),
    .C1(_0948_),
    .D1(_0950_),
    .X(_0951_)
  );
  sky130_fd_sc_hd__and3_2 _3274_ (
    .A(\g_bit[10].g_word[27].r_bit.Q ),
    .B(_0852_),
    .C(_0853_),
    .X(_0952_)
  );
  sky130_fd_sc_hd__a221o_2 _3275_ (
    .A1(\g_bit[10].g_word[6].r_bit.Q ),
    .A2(_0850_),
    .B1(_0851_),
    .B2(\g_bit[10].g_word[1].r_bit.Q ),
    .C1(_0952_),
    .X(_0953_)
  );
  sky130_fd_sc_hd__inv_2 _3276_ (
    .A(\g_bit[10].g_word[23].r_bit.Q ),
    .Y(_0954_)
  );
  sky130_fd_sc_hd__inv_2 _3277_ (
    .A(\g_bit[10].g_word[10].r_bit.Q ),
    .Y(_0955_)
  );
  sky130_fd_sc_hd__or3_2 _3278_ (
    .A(_0955_),
    .B(_0453_),
    .C(_0700_),
    .X(_0956_)
  );
  sky130_fd_sc_hd__inv_2 _3279_ (
    .A(\g_bit[10].g_word[9].r_bit.Q ),
    .Y(_0957_)
  );
  sky130_fd_sc_hd__or3_2 _3280_ (
    .A(_0957_),
    .B(_0577_),
    .C(_0861_),
    .X(_0958_)
  );
  sky130_fd_sc_hd__inv_2 _3281_ (
    .A(\g_bit[10].g_word[8].r_bit.Q ),
    .Y(_0959_)
  );
  sky130_fd_sc_hd__or3_2 _3282_ (
    .A(_0959_),
    .B(_0705_),
    .C(_0864_),
    .X(_0960_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3283_ (
    .A1(_0954_),
    .A2(_0857_),
    .B1(_0956_),
    .C1(_0958_),
    .D1(_0960_),
    .Y(_0961_)
  );
  sky130_fd_sc_hd__inv_2 _3284_ (
    .A(\g_bit[10].g_word[22].r_bit.Q ),
    .Y(_0962_)
  );
  sky130_fd_sc_hd__inv_2 _3285_ (
    .A(\g_bit[10].g_word[16].r_bit.Q ),
    .Y(_0963_)
  );
  sky130_fd_sc_hd__or3_2 _3286_ (
    .A(_0963_),
    .B(_0584_),
    .C(_0870_),
    .X(_0964_)
  );
  sky130_fd_sc_hd__inv_2 _3287_ (
    .A(\g_bit[10].g_word[14].r_bit.Q ),
    .Y(_0965_)
  );
  sky130_fd_sc_hd__or3_2 _3288_ (
    .A(_0965_),
    .B(_0873_),
    .C(_0777_),
    .X(_0966_)
  );
  sky130_fd_sc_hd__inv_2 _3289_ (
    .A(\g_bit[10].g_word[18].r_bit.Q ),
    .Y(_0967_)
  );
  sky130_fd_sc_hd__or3_2 _3290_ (
    .A(_0967_),
    .B(_0780_),
    .C(_0876_),
    .X(_0968_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3291_ (
    .A1(_0962_),
    .A2(_0868_),
    .B1(_0964_),
    .C1(_0966_),
    .D1(_0968_),
    .Y(_0969_)
  );
  sky130_fd_sc_hd__or4_2 _3292_ (
    .A(_0951_),
    .B(_0953_),
    .C(_0961_),
    .D(_0969_),
    .X(_0970_)
  );
  sky130_fd_sc_hd__or4_2 _3293_ (
    .A(_0937_),
    .B(_0939_),
    .C(_0944_),
    .D(_0970_),
    .X(_0971_)
  );
  sky130_fd_sc_hd__buf_1 _3294_ (
    .A(_0971_),
    .X(\g_bit[10].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _3295_ (
    .A1(\g_bit[10].g_word[30].r_bit.Q ),
    .A2(_0883_),
    .A3(_0884_),
    .B1(_0885_),
    .B2(\g_bit[10].g_word[28].r_bit.Q ),
    .X(_0972_)
  );
  sky130_fd_sc_hd__a221o_2 _3296_ (
    .A1(\g_bit[10].g_word[4].r_bit.Q ),
    .A2(_0881_),
    .B1(_0882_),
    .B2(\g_bit[10].g_word[26].r_bit.Q ),
    .C1(_0972_),
    .X(_0973_)
  );
  sky130_fd_sc_hd__a22o_2 _3297_ (
    .A1(\g_bit[10].g_word[5].r_bit.Q ),
    .A2(_0890_),
    .B1(_0891_),
    .B2(\g_bit[10].g_word[2].r_bit.Q ),
    .X(_0974_)
  );
  sky130_fd_sc_hd__a221o_2 _3298_ (
    .A1(\g_bit[10].g_word[25].r_bit.Q ),
    .A2(_0888_),
    .B1(_0889_),
    .B2(\g_bit[10].g_word[31].r_bit.Q ),
    .C1(_0974_),
    .X(_0975_)
  );
  sky130_fd_sc_hd__a22o_2 _3299_ (
    .A1(\g_bit[10].g_word[13].r_bit.Q ),
    .A2(_0894_),
    .B1(_0895_),
    .B2(\g_bit[10].g_word[15].r_bit.Q ),
    .X(_0976_)
  );
  sky130_fd_sc_hd__a22o_2 _3300_ (
    .A1(\g_bit[10].g_word[20].r_bit.Q ),
    .A2(_0897_),
    .B1(_0898_),
    .B2(\g_bit[10].g_word[11].r_bit.Q ),
    .X(_0977_)
  );
  sky130_fd_sc_hd__a22o_2 _3301_ (
    .A1(\g_bit[10].g_word[19].r_bit.Q ),
    .A2(_0900_),
    .B1(_0901_),
    .B2(\g_bit[10].g_word[21].r_bit.Q ),
    .X(_0978_)
  );
  sky130_fd_sc_hd__a22o_2 _3302_ (
    .A1(\g_bit[10].g_word[17].r_bit.Q ),
    .A2(_0903_),
    .B1(_0904_),
    .B2(\g_bit[10].g_word[12].r_bit.Q ),
    .X(_0979_)
  );
  sky130_fd_sc_hd__or4_2 _3303_ (
    .A(_0976_),
    .B(_0977_),
    .C(_0978_),
    .D(_0979_),
    .X(_0980_)
  );
  sky130_fd_sc_hd__nor3_2 _3304_ (
    .A(_0945_),
    .B(_0794_),
    .C(_0727_),
    .Y(_0981_)
  );
  sky130_fd_sc_hd__nor3_2 _3305_ (
    .A(_0947_),
    .B(_0909_),
    .C(_0796_),
    .Y(_0982_)
  );
  sky130_fd_sc_hd__buf_1 _3306_ (
    .A(_0206_),
    .X(_0983_)
  );
  sky130_fd_sc_hd__and3_2 _3307_ (
    .A(\g_bit[10].g_word[24].r_bit.Q ),
    .B(_0983_),
    .C(_0798_),
    .X(_0984_)
  );
  sky130_fd_sc_hd__a2111o_2 _3308_ (
    .A1(\g_bit[10].g_word[29].r_bit.Q ),
    .A2(_0907_),
    .B1(_0981_),
    .C1(_0982_),
    .D1(_0984_),
    .X(_0985_)
  );
  sky130_fd_sc_hd__and3_2 _3309_ (
    .A(\g_bit[10].g_word[27].r_bit.Q ),
    .B(_0915_),
    .C(_0916_),
    .X(_0986_)
  );
  sky130_fd_sc_hd__a221o_2 _3310_ (
    .A1(\g_bit[10].g_word[6].r_bit.Q ),
    .A2(_0913_),
    .B1(_0914_),
    .B2(\g_bit[10].g_word[1].r_bit.Q ),
    .C1(_0986_),
    .X(_0987_)
  );
  sky130_fd_sc_hd__or3_2 _3311_ (
    .A(_0955_),
    .B(_0485_),
    .C(_0734_),
    .X(_0988_)
  );
  sky130_fd_sc_hd__or3_2 _3312_ (
    .A(_0957_),
    .B(_0609_),
    .C(_0921_),
    .X(_0989_)
  );
  sky130_fd_sc_hd__or3_2 _3313_ (
    .A(_0959_),
    .B(_0737_),
    .C(_0923_),
    .X(_0990_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3314_ (
    .A1(_0954_),
    .A2(_0919_),
    .B1(_0988_),
    .C1(_0989_),
    .D1(_0990_),
    .Y(_0991_)
  );
  sky130_fd_sc_hd__or3_2 _3315_ (
    .A(_0963_),
    .B(_0927_),
    .C(_0673_),
    .X(_0992_)
  );
  sky130_fd_sc_hd__or3_2 _3316_ (
    .A(_0965_),
    .B(_0929_),
    .C(_0808_),
    .X(_0993_)
  );
  sky130_fd_sc_hd__or3_2 _3317_ (
    .A(_0967_),
    .B(_0810_),
    .C(_0931_),
    .X(_0994_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3318_ (
    .A1(_0962_),
    .A2(_0926_),
    .B1(_0992_),
    .C1(_0993_),
    .D1(_0994_),
    .Y(_0995_)
  );
  sky130_fd_sc_hd__or4_2 _3319_ (
    .A(_0985_),
    .B(_0987_),
    .C(_0991_),
    .D(_0995_),
    .X(_0996_)
  );
  sky130_fd_sc_hd__or4_2 _3320_ (
    .A(_0973_),
    .B(_0975_),
    .C(_0980_),
    .D(_0996_),
    .X(_0997_)
  );
  sky130_fd_sc_hd__buf_1 _3321_ (
    .A(_0997_),
    .X(\g_bit[10].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _3322_ (
    .A1(\g_bit[11].g_word[30].r_bit.Q ),
    .A2(_0817_),
    .A3(_0818_),
    .B1(_0819_),
    .B2(\g_bit[11].g_word[28].r_bit.Q ),
    .X(_0998_)
  );
  sky130_fd_sc_hd__a221o_2 _3323_ (
    .A1(\g_bit[11].g_word[4].r_bit.Q ),
    .A2(_0815_),
    .B1(_0816_),
    .B2(\g_bit[11].g_word[26].r_bit.Q ),
    .C1(_0998_),
    .X(_0999_)
  );
  sky130_fd_sc_hd__a22o_2 _3324_ (
    .A1(\g_bit[11].g_word[5].r_bit.Q ),
    .A2(_0824_),
    .B1(_0825_),
    .B2(\g_bit[11].g_word[2].r_bit.Q ),
    .X(_1000_)
  );
  sky130_fd_sc_hd__a221o_2 _3325_ (
    .A1(\g_bit[11].g_word[25].r_bit.Q ),
    .A2(_0822_),
    .B1(_0823_),
    .B2(\g_bit[11].g_word[31].r_bit.Q ),
    .C1(_1000_),
    .X(_1001_)
  );
  sky130_fd_sc_hd__a22o_2 _3326_ (
    .A1(\g_bit[11].g_word[13].r_bit.Q ),
    .A2(_0828_),
    .B1(_0829_),
    .B2(\g_bit[11].g_word[15].r_bit.Q ),
    .X(_1002_)
  );
  sky130_fd_sc_hd__a22o_2 _3327_ (
    .A1(\g_bit[11].g_word[11].r_bit.Q ),
    .A2(_0831_),
    .B1(_0832_),
    .B2(\g_bit[11].g_word[20].r_bit.Q ),
    .X(_1003_)
  );
  sky130_fd_sc_hd__a22o_2 _3328_ (
    .A1(\g_bit[11].g_word[19].r_bit.Q ),
    .A2(_0834_),
    .B1(_0835_),
    .B2(\g_bit[11].g_word[21].r_bit.Q ),
    .X(_1004_)
  );
  sky130_fd_sc_hd__a22o_2 _3329_ (
    .A1(\g_bit[11].g_word[17].r_bit.Q ),
    .A2(_0837_),
    .B1(_0838_),
    .B2(\g_bit[11].g_word[12].r_bit.Q ),
    .X(_1005_)
  );
  sky130_fd_sc_hd__or4_2 _3330_ (
    .A(_1002_),
    .B(_1003_),
    .C(_1004_),
    .D(_1005_),
    .X(_1006_)
  );
  sky130_fd_sc_hd__inv_2 _3331_ (
    .A(\g_bit[11].g_word[7].r_bit.Q ),
    .Y(_1007_)
  );
  sky130_fd_sc_hd__nor3_2 _3332_ (
    .A(_1007_),
    .B(_0690_),
    .C(_0756_),
    .Y(_1008_)
  );
  sky130_fd_sc_hd__inv_2 _3333_ (
    .A(\g_bit[11].g_word[3].r_bit.Q ),
    .Y(_1009_)
  );
  sky130_fd_sc_hd__nor3_2 _3334_ (
    .A(_1009_),
    .B(_0845_),
    .C(_0846_),
    .Y(_1010_)
  );
  sky130_fd_sc_hd__and3_2 _3335_ (
    .A(\g_bit[11].g_word[24].r_bit.Q ),
    .B(_0760_),
    .C(_0949_),
    .X(_1011_)
  );
  sky130_fd_sc_hd__a2111o_2 _3336_ (
    .A1(\g_bit[11].g_word[29].r_bit.Q ),
    .A2(_0841_),
    .B1(_1008_),
    .C1(_1010_),
    .D1(_1011_),
    .X(_1012_)
  );
  sky130_fd_sc_hd__and3_2 _3337_ (
    .A(\g_bit[11].g_word[27].r_bit.Q ),
    .B(_0852_),
    .C(_0853_),
    .X(_1013_)
  );
  sky130_fd_sc_hd__a221o_2 _3338_ (
    .A1(\g_bit[11].g_word[6].r_bit.Q ),
    .A2(_0850_),
    .B1(_0851_),
    .B2(\g_bit[11].g_word[1].r_bit.Q ),
    .C1(_1013_),
    .X(_1014_)
  );
  sky130_fd_sc_hd__inv_2 _3339_ (
    .A(\g_bit[11].g_word[23].r_bit.Q ),
    .Y(_1015_)
  );
  sky130_fd_sc_hd__inv_2 _3340_ (
    .A(\g_bit[11].g_word[10].r_bit.Q ),
    .Y(_1016_)
  );
  sky130_fd_sc_hd__or3_2 _3341_ (
    .A(_1016_),
    .B(_0453_),
    .C(_0700_),
    .X(_1017_)
  );
  sky130_fd_sc_hd__inv_2 _3342_ (
    .A(\g_bit[11].g_word[9].r_bit.Q ),
    .Y(_1018_)
  );
  sky130_fd_sc_hd__or3_2 _3343_ (
    .A(_1018_),
    .B(_0577_),
    .C(_0861_),
    .X(_1019_)
  );
  sky130_fd_sc_hd__inv_2 _3344_ (
    .A(\g_bit[11].g_word[8].r_bit.Q ),
    .Y(_1020_)
  );
  sky130_fd_sc_hd__or3_2 _3345_ (
    .A(_1020_),
    .B(_0705_),
    .C(_0864_),
    .X(_1021_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3346_ (
    .A1(_1015_),
    .A2(_0857_),
    .B1(_1017_),
    .C1(_1019_),
    .D1(_1021_),
    .Y(_1022_)
  );
  sky130_fd_sc_hd__inv_2 _3347_ (
    .A(\g_bit[11].g_word[22].r_bit.Q ),
    .Y(_1023_)
  );
  sky130_fd_sc_hd__inv_2 _3348_ (
    .A(\g_bit[11].g_word[16].r_bit.Q ),
    .Y(_1024_)
  );
  sky130_fd_sc_hd__or3_2 _3349_ (
    .A(_1024_),
    .B(_0584_),
    .C(_0870_),
    .X(_1025_)
  );
  sky130_fd_sc_hd__inv_2 _3350_ (
    .A(\g_bit[11].g_word[14].r_bit.Q ),
    .Y(_1026_)
  );
  sky130_fd_sc_hd__or3_2 _3351_ (
    .A(_1026_),
    .B(_0873_),
    .C(_0777_),
    .X(_1027_)
  );
  sky130_fd_sc_hd__inv_2 _3352_ (
    .A(\g_bit[11].g_word[18].r_bit.Q ),
    .Y(_1028_)
  );
  sky130_fd_sc_hd__or3_2 _3353_ (
    .A(_1028_),
    .B(_0780_),
    .C(_0876_),
    .X(_1029_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3354_ (
    .A1(_1023_),
    .A2(_0868_),
    .B1(_1025_),
    .C1(_1027_),
    .D1(_1029_),
    .Y(_1030_)
  );
  sky130_fd_sc_hd__or4_2 _3355_ (
    .A(_1012_),
    .B(_1014_),
    .C(_1022_),
    .D(_1030_),
    .X(_1031_)
  );
  sky130_fd_sc_hd__or4_2 _3356_ (
    .A(_0999_),
    .B(_1001_),
    .C(_1006_),
    .D(_1031_),
    .X(_1032_)
  );
  sky130_fd_sc_hd__buf_1 _3357_ (
    .A(_1032_),
    .X(\g_bit[11].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _3358_ (
    .A1(\g_bit[11].g_word[30].r_bit.Q ),
    .A2(_0883_),
    .A3(_0884_),
    .B1(_0885_),
    .B2(\g_bit[11].g_word[28].r_bit.Q ),
    .X(_1033_)
  );
  sky130_fd_sc_hd__a221o_2 _3359_ (
    .A1(\g_bit[11].g_word[4].r_bit.Q ),
    .A2(_0881_),
    .B1(_0882_),
    .B2(\g_bit[11].g_word[26].r_bit.Q ),
    .C1(_1033_),
    .X(_1034_)
  );
  sky130_fd_sc_hd__a22o_2 _3360_ (
    .A1(\g_bit[11].g_word[5].r_bit.Q ),
    .A2(_0890_),
    .B1(_0891_),
    .B2(\g_bit[11].g_word[2].r_bit.Q ),
    .X(_1035_)
  );
  sky130_fd_sc_hd__a221o_2 _3361_ (
    .A1(\g_bit[11].g_word[25].r_bit.Q ),
    .A2(_0888_),
    .B1(_0889_),
    .B2(\g_bit[11].g_word[31].r_bit.Q ),
    .C1(_1035_),
    .X(_1036_)
  );
  sky130_fd_sc_hd__a22o_2 _3362_ (
    .A1(\g_bit[11].g_word[13].r_bit.Q ),
    .A2(_0894_),
    .B1(_0895_),
    .B2(\g_bit[11].g_word[15].r_bit.Q ),
    .X(_1037_)
  );
  sky130_fd_sc_hd__a22o_2 _3363_ (
    .A1(\g_bit[11].g_word[20].r_bit.Q ),
    .A2(_0897_),
    .B1(_0898_),
    .B2(\g_bit[11].g_word[11].r_bit.Q ),
    .X(_1038_)
  );
  sky130_fd_sc_hd__a22o_2 _3364_ (
    .A1(\g_bit[11].g_word[19].r_bit.Q ),
    .A2(_0900_),
    .B1(_0901_),
    .B2(\g_bit[11].g_word[21].r_bit.Q ),
    .X(_1039_)
  );
  sky130_fd_sc_hd__a22o_2 _3365_ (
    .A1(\g_bit[11].g_word[17].r_bit.Q ),
    .A2(_0903_),
    .B1(_0904_),
    .B2(\g_bit[11].g_word[12].r_bit.Q ),
    .X(_1040_)
  );
  sky130_fd_sc_hd__or4_2 _3366_ (
    .A(_1037_),
    .B(_1038_),
    .C(_1039_),
    .D(_1040_),
    .X(_1041_)
  );
  sky130_fd_sc_hd__nor3_2 _3367_ (
    .A(_1007_),
    .B(_0794_),
    .C(_0727_),
    .Y(_1042_)
  );
  sky130_fd_sc_hd__nor3_2 _3368_ (
    .A(_1009_),
    .B(_0909_),
    .C(_0796_),
    .Y(_1043_)
  );
  sky130_fd_sc_hd__and3_2 _3369_ (
    .A(\g_bit[11].g_word[24].r_bit.Q ),
    .B(_0983_),
    .C(_0798_),
    .X(_1044_)
  );
  sky130_fd_sc_hd__a2111o_2 _3370_ (
    .A1(\g_bit[11].g_word[29].r_bit.Q ),
    .A2(_0907_),
    .B1(_1042_),
    .C1(_1043_),
    .D1(_1044_),
    .X(_1045_)
  );
  sky130_fd_sc_hd__and3_2 _3371_ (
    .A(\g_bit[11].g_word[27].r_bit.Q ),
    .B(_0915_),
    .C(_0916_),
    .X(_1046_)
  );
  sky130_fd_sc_hd__a221o_2 _3372_ (
    .A1(\g_bit[11].g_word[6].r_bit.Q ),
    .A2(_0913_),
    .B1(_0914_),
    .B2(\g_bit[11].g_word[1].r_bit.Q ),
    .C1(_1046_),
    .X(_1047_)
  );
  sky130_fd_sc_hd__or3_2 _3373_ (
    .A(_1016_),
    .B(_0485_),
    .C(_0734_),
    .X(_1048_)
  );
  sky130_fd_sc_hd__or3_2 _3374_ (
    .A(_1018_),
    .B(_0609_),
    .C(_0921_),
    .X(_1049_)
  );
  sky130_fd_sc_hd__or3_2 _3375_ (
    .A(_1020_),
    .B(_0737_),
    .C(_0923_),
    .X(_1050_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3376_ (
    .A1(_1015_),
    .A2(_0919_),
    .B1(_1048_),
    .C1(_1049_),
    .D1(_1050_),
    .Y(_1051_)
  );
  sky130_fd_sc_hd__or3_2 _3377_ (
    .A(_1024_),
    .B(_0927_),
    .C(_0673_),
    .X(_1052_)
  );
  sky130_fd_sc_hd__or3_2 _3378_ (
    .A(_1026_),
    .B(_0929_),
    .C(_0808_),
    .X(_1053_)
  );
  sky130_fd_sc_hd__or3_2 _3379_ (
    .A(_1028_),
    .B(_0810_),
    .C(_0931_),
    .X(_1054_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3380_ (
    .A1(_1023_),
    .A2(_0926_),
    .B1(_1052_),
    .C1(_1053_),
    .D1(_1054_),
    .Y(_1055_)
  );
  sky130_fd_sc_hd__or4_2 _3381_ (
    .A(_1045_),
    .B(_1047_),
    .C(_1051_),
    .D(_1055_),
    .X(_1056_)
  );
  sky130_fd_sc_hd__or4_2 _3382_ (
    .A(_1034_),
    .B(_1036_),
    .C(_1041_),
    .D(_1056_),
    .X(_1057_)
  );
  sky130_fd_sc_hd__buf_1 _3383_ (
    .A(_1057_),
    .X(\g_bit[11].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _3384_ (
    .A1(\g_bit[12].g_word[30].r_bit.Q ),
    .A2(_0817_),
    .A3(_0818_),
    .B1(_0819_),
    .B2(\g_bit[12].g_word[28].r_bit.Q ),
    .X(_1058_)
  );
  sky130_fd_sc_hd__a221o_2 _3385_ (
    .A1(\g_bit[12].g_word[4].r_bit.Q ),
    .A2(_0815_),
    .B1(_0816_),
    .B2(\g_bit[12].g_word[26].r_bit.Q ),
    .C1(_1058_),
    .X(_1059_)
  );
  sky130_fd_sc_hd__a22o_2 _3386_ (
    .A1(\g_bit[12].g_word[5].r_bit.Q ),
    .A2(_0824_),
    .B1(_0825_),
    .B2(\g_bit[12].g_word[2].r_bit.Q ),
    .X(_1060_)
  );
  sky130_fd_sc_hd__a221o_2 _3387_ (
    .A1(\g_bit[12].g_word[25].r_bit.Q ),
    .A2(_0822_),
    .B1(_0823_),
    .B2(\g_bit[12].g_word[31].r_bit.Q ),
    .C1(_1060_),
    .X(_1061_)
  );
  sky130_fd_sc_hd__a22o_2 _3388_ (
    .A1(\g_bit[12].g_word[13].r_bit.Q ),
    .A2(_0828_),
    .B1(_0829_),
    .B2(\g_bit[12].g_word[15].r_bit.Q ),
    .X(_1062_)
  );
  sky130_fd_sc_hd__a22o_2 _3389_ (
    .A1(\g_bit[12].g_word[11].r_bit.Q ),
    .A2(_0831_),
    .B1(_0832_),
    .B2(\g_bit[12].g_word[20].r_bit.Q ),
    .X(_1063_)
  );
  sky130_fd_sc_hd__a22o_2 _3390_ (
    .A1(\g_bit[12].g_word[19].r_bit.Q ),
    .A2(_0834_),
    .B1(_0835_),
    .B2(\g_bit[12].g_word[21].r_bit.Q ),
    .X(_1064_)
  );
  sky130_fd_sc_hd__a22o_2 _3391_ (
    .A1(\g_bit[12].g_word[17].r_bit.Q ),
    .A2(_0837_),
    .B1(_0838_),
    .B2(\g_bit[12].g_word[12].r_bit.Q ),
    .X(_1065_)
  );
  sky130_fd_sc_hd__or4_2 _3392_ (
    .A(_1062_),
    .B(_1063_),
    .C(_1064_),
    .D(_1065_),
    .X(_1066_)
  );
  sky130_fd_sc_hd__inv_2 _3393_ (
    .A(\g_bit[12].g_word[7].r_bit.Q ),
    .Y(_1067_)
  );
  sky130_fd_sc_hd__nor3_2 _3394_ (
    .A(_1067_),
    .B(_0690_),
    .C(_0756_),
    .Y(_1068_)
  );
  sky130_fd_sc_hd__inv_2 _3395_ (
    .A(\g_bit[12].g_word[3].r_bit.Q ),
    .Y(_1069_)
  );
  sky130_fd_sc_hd__nor3_2 _3396_ (
    .A(_1069_),
    .B(_0845_),
    .C(_0846_),
    .Y(_1070_)
  );
  sky130_fd_sc_hd__and3_2 _3397_ (
    .A(\g_bit[12].g_word[24].r_bit.Q ),
    .B(_0760_),
    .C(_0949_),
    .X(_1071_)
  );
  sky130_fd_sc_hd__a2111o_2 _3398_ (
    .A1(\g_bit[12].g_word[29].r_bit.Q ),
    .A2(_0841_),
    .B1(_1068_),
    .C1(_1070_),
    .D1(_1071_),
    .X(_1072_)
  );
  sky130_fd_sc_hd__and3_2 _3399_ (
    .A(\g_bit[12].g_word[27].r_bit.Q ),
    .B(_0852_),
    .C(_0853_),
    .X(_1073_)
  );
  sky130_fd_sc_hd__a221o_2 _3400_ (
    .A1(\g_bit[12].g_word[6].r_bit.Q ),
    .A2(_0850_),
    .B1(_0851_),
    .B2(\g_bit[12].g_word[1].r_bit.Q ),
    .C1(_1073_),
    .X(_1074_)
  );
  sky130_fd_sc_hd__inv_2 _3401_ (
    .A(\g_bit[12].g_word[23].r_bit.Q ),
    .Y(_1075_)
  );
  sky130_fd_sc_hd__inv_2 _3402_ (
    .A(\g_bit[12].g_word[10].r_bit.Q ),
    .Y(_1076_)
  );
  sky130_fd_sc_hd__or3_2 _3403_ (
    .A(_1076_),
    .B(_0453_),
    .C(_0700_),
    .X(_1077_)
  );
  sky130_fd_sc_hd__inv_2 _3404_ (
    .A(\g_bit[12].g_word[9].r_bit.Q ),
    .Y(_1078_)
  );
  sky130_fd_sc_hd__or3_2 _3405_ (
    .A(_1078_),
    .B(_0577_),
    .C(_0861_),
    .X(_1079_)
  );
  sky130_fd_sc_hd__inv_2 _3406_ (
    .A(\g_bit[12].g_word[8].r_bit.Q ),
    .Y(_1080_)
  );
  sky130_fd_sc_hd__or3_2 _3407_ (
    .A(_1080_),
    .B(_0705_),
    .C(_0864_),
    .X(_1081_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3408_ (
    .A1(_1075_),
    .A2(_0857_),
    .B1(_1077_),
    .C1(_1079_),
    .D1(_1081_),
    .Y(_1082_)
  );
  sky130_fd_sc_hd__inv_2 _3409_ (
    .A(\g_bit[12].g_word[22].r_bit.Q ),
    .Y(_1083_)
  );
  sky130_fd_sc_hd__inv_2 _3410_ (
    .A(\g_bit[12].g_word[16].r_bit.Q ),
    .Y(_1084_)
  );
  sky130_fd_sc_hd__or3_2 _3411_ (
    .A(_1084_),
    .B(_0584_),
    .C(_0870_),
    .X(_1085_)
  );
  sky130_fd_sc_hd__inv_2 _3412_ (
    .A(\g_bit[12].g_word[14].r_bit.Q ),
    .Y(_1086_)
  );
  sky130_fd_sc_hd__or3_2 _3413_ (
    .A(_1086_),
    .B(_0873_),
    .C(_0777_),
    .X(_1087_)
  );
  sky130_fd_sc_hd__inv_2 _3414_ (
    .A(\g_bit[12].g_word[18].r_bit.Q ),
    .Y(_1088_)
  );
  sky130_fd_sc_hd__or3_2 _3415_ (
    .A(_1088_),
    .B(_0780_),
    .C(_0876_),
    .X(_1089_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3416_ (
    .A1(_1083_),
    .A2(_0868_),
    .B1(_1085_),
    .C1(_1087_),
    .D1(_1089_),
    .Y(_1090_)
  );
  sky130_fd_sc_hd__or4_2 _3417_ (
    .A(_1072_),
    .B(_1074_),
    .C(_1082_),
    .D(_1090_),
    .X(_1091_)
  );
  sky130_fd_sc_hd__or4_2 _3418_ (
    .A(_1059_),
    .B(_1061_),
    .C(_1066_),
    .D(_1091_),
    .X(_1092_)
  );
  sky130_fd_sc_hd__buf_1 _3419_ (
    .A(_1092_),
    .X(\g_bit[12].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _3420_ (
    .A1(\g_bit[12].g_word[30].r_bit.Q ),
    .A2(_0883_),
    .A3(_0884_),
    .B1(_0885_),
    .B2(\g_bit[12].g_word[28].r_bit.Q ),
    .X(_1093_)
  );
  sky130_fd_sc_hd__a221o_2 _3421_ (
    .A1(\g_bit[12].g_word[4].r_bit.Q ),
    .A2(_0881_),
    .B1(_0882_),
    .B2(\g_bit[12].g_word[26].r_bit.Q ),
    .C1(_1093_),
    .X(_1094_)
  );
  sky130_fd_sc_hd__a22o_2 _3422_ (
    .A1(\g_bit[12].g_word[5].r_bit.Q ),
    .A2(_0890_),
    .B1(_0891_),
    .B2(\g_bit[12].g_word[2].r_bit.Q ),
    .X(_1095_)
  );
  sky130_fd_sc_hd__a221o_2 _3423_ (
    .A1(\g_bit[12].g_word[25].r_bit.Q ),
    .A2(_0888_),
    .B1(_0889_),
    .B2(\g_bit[12].g_word[31].r_bit.Q ),
    .C1(_1095_),
    .X(_1096_)
  );
  sky130_fd_sc_hd__a22o_2 _3424_ (
    .A1(\g_bit[12].g_word[13].r_bit.Q ),
    .A2(_0894_),
    .B1(_0895_),
    .B2(\g_bit[12].g_word[15].r_bit.Q ),
    .X(_1097_)
  );
  sky130_fd_sc_hd__a22o_2 _3425_ (
    .A1(\g_bit[12].g_word[20].r_bit.Q ),
    .A2(_0897_),
    .B1(_0898_),
    .B2(\g_bit[12].g_word[11].r_bit.Q ),
    .X(_1098_)
  );
  sky130_fd_sc_hd__a22o_2 _3426_ (
    .A1(\g_bit[12].g_word[19].r_bit.Q ),
    .A2(_0900_),
    .B1(_0901_),
    .B2(\g_bit[12].g_word[21].r_bit.Q ),
    .X(_1099_)
  );
  sky130_fd_sc_hd__a22o_2 _3427_ (
    .A1(\g_bit[12].g_word[17].r_bit.Q ),
    .A2(_0903_),
    .B1(_0904_),
    .B2(\g_bit[12].g_word[12].r_bit.Q ),
    .X(_1100_)
  );
  sky130_fd_sc_hd__or4_2 _3428_ (
    .A(_1097_),
    .B(_1098_),
    .C(_1099_),
    .D(_1100_),
    .X(_1101_)
  );
  sky130_fd_sc_hd__nor3_2 _3429_ (
    .A(_1067_),
    .B(_0794_),
    .C(_0727_),
    .Y(_1102_)
  );
  sky130_fd_sc_hd__nor3_2 _3430_ (
    .A(_1069_),
    .B(_0909_),
    .C(_0796_),
    .Y(_1103_)
  );
  sky130_fd_sc_hd__and3_2 _3431_ (
    .A(\g_bit[12].g_word[24].r_bit.Q ),
    .B(_0983_),
    .C(_0798_),
    .X(_1104_)
  );
  sky130_fd_sc_hd__a2111o_2 _3432_ (
    .A1(\g_bit[12].g_word[29].r_bit.Q ),
    .A2(_0907_),
    .B1(_1102_),
    .C1(_1103_),
    .D1(_1104_),
    .X(_1105_)
  );
  sky130_fd_sc_hd__and3_2 _3433_ (
    .A(\g_bit[12].g_word[27].r_bit.Q ),
    .B(_0915_),
    .C(_0916_),
    .X(_1106_)
  );
  sky130_fd_sc_hd__a221o_2 _3434_ (
    .A1(\g_bit[12].g_word[6].r_bit.Q ),
    .A2(_0913_),
    .B1(_0914_),
    .B2(\g_bit[12].g_word[1].r_bit.Q ),
    .C1(_1106_),
    .X(_1107_)
  );
  sky130_fd_sc_hd__or3_2 _3435_ (
    .A(_1076_),
    .B(_0485_),
    .C(_0734_),
    .X(_1108_)
  );
  sky130_fd_sc_hd__or3_2 _3436_ (
    .A(_1078_),
    .B(_0609_),
    .C(_0921_),
    .X(_1109_)
  );
  sky130_fd_sc_hd__or3_2 _3437_ (
    .A(_1080_),
    .B(_0737_),
    .C(_0923_),
    .X(_1110_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3438_ (
    .A1(_1075_),
    .A2(_0919_),
    .B1(_1108_),
    .C1(_1109_),
    .D1(_1110_),
    .Y(_1111_)
  );
  sky130_fd_sc_hd__or3_2 _3439_ (
    .A(_1084_),
    .B(_0927_),
    .C(_0673_),
    .X(_1112_)
  );
  sky130_fd_sc_hd__or3_2 _3440_ (
    .A(_1086_),
    .B(_0929_),
    .C(_0808_),
    .X(_1113_)
  );
  sky130_fd_sc_hd__or3_2 _3441_ (
    .A(_1088_),
    .B(_0810_),
    .C(_0931_),
    .X(_1114_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3442_ (
    .A1(_1083_),
    .A2(_0926_),
    .B1(_1112_),
    .C1(_1113_),
    .D1(_1114_),
    .Y(_1115_)
  );
  sky130_fd_sc_hd__or4_2 _3443_ (
    .A(_1105_),
    .B(_1107_),
    .C(_1111_),
    .D(_1115_),
    .X(_1116_)
  );
  sky130_fd_sc_hd__or4_2 _3444_ (
    .A(_1094_),
    .B(_1096_),
    .C(_1101_),
    .D(_1116_),
    .X(_1117_)
  );
  sky130_fd_sc_hd__buf_1 _3445_ (
    .A(_1117_),
    .X(\g_bit[12].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _3446_ (
    .A1(\g_bit[13].g_word[30].r_bit.Q ),
    .A2(_0817_),
    .A3(_0818_),
    .B1(_0819_),
    .B2(\g_bit[13].g_word[28].r_bit.Q ),
    .X(_1118_)
  );
  sky130_fd_sc_hd__a221o_2 _3447_ (
    .A1(\g_bit[13].g_word[4].r_bit.Q ),
    .A2(_0815_),
    .B1(_0816_),
    .B2(\g_bit[13].g_word[26].r_bit.Q ),
    .C1(_1118_),
    .X(_1119_)
  );
  sky130_fd_sc_hd__a22o_2 _3448_ (
    .A1(\g_bit[13].g_word[5].r_bit.Q ),
    .A2(_0824_),
    .B1(_0825_),
    .B2(\g_bit[13].g_word[2].r_bit.Q ),
    .X(_1120_)
  );
  sky130_fd_sc_hd__a221o_2 _3449_ (
    .A1(\g_bit[13].g_word[25].r_bit.Q ),
    .A2(_0822_),
    .B1(_0823_),
    .B2(\g_bit[13].g_word[31].r_bit.Q ),
    .C1(_1120_),
    .X(_1121_)
  );
  sky130_fd_sc_hd__a22o_2 _3450_ (
    .A1(\g_bit[13].g_word[13].r_bit.Q ),
    .A2(_0828_),
    .B1(_0829_),
    .B2(\g_bit[13].g_word[15].r_bit.Q ),
    .X(_1122_)
  );
  sky130_fd_sc_hd__a22o_2 _3451_ (
    .A1(\g_bit[13].g_word[11].r_bit.Q ),
    .A2(_0831_),
    .B1(_0832_),
    .B2(\g_bit[13].g_word[20].r_bit.Q ),
    .X(_1123_)
  );
  sky130_fd_sc_hd__a22o_2 _3452_ (
    .A1(\g_bit[13].g_word[19].r_bit.Q ),
    .A2(_0834_),
    .B1(_0835_),
    .B2(\g_bit[13].g_word[21].r_bit.Q ),
    .X(_1124_)
  );
  sky130_fd_sc_hd__a22o_2 _3453_ (
    .A1(\g_bit[13].g_word[17].r_bit.Q ),
    .A2(_0837_),
    .B1(_0838_),
    .B2(\g_bit[13].g_word[12].r_bit.Q ),
    .X(_1125_)
  );
  sky130_fd_sc_hd__or4_2 _3454_ (
    .A(_1122_),
    .B(_1123_),
    .C(_1124_),
    .D(_1125_),
    .X(_1126_)
  );
  sky130_fd_sc_hd__inv_2 _3455_ (
    .A(\g_bit[13].g_word[7].r_bit.Q ),
    .Y(_1127_)
  );
  sky130_fd_sc_hd__nor3_2 _3456_ (
    .A(_1127_),
    .B(_0690_),
    .C(_0756_),
    .Y(_1128_)
  );
  sky130_fd_sc_hd__inv_2 _3457_ (
    .A(\g_bit[13].g_word[3].r_bit.Q ),
    .Y(_1129_)
  );
  sky130_fd_sc_hd__nor3_2 _3458_ (
    .A(_1129_),
    .B(_0845_),
    .C(_0846_),
    .Y(_1130_)
  );
  sky130_fd_sc_hd__and3_2 _3459_ (
    .A(\g_bit[13].g_word[24].r_bit.Q ),
    .B(_0760_),
    .C(_0949_),
    .X(_1131_)
  );
  sky130_fd_sc_hd__a2111o_2 _3460_ (
    .A1(\g_bit[13].g_word[29].r_bit.Q ),
    .A2(_0841_),
    .B1(_1128_),
    .C1(_1130_),
    .D1(_1131_),
    .X(_1132_)
  );
  sky130_fd_sc_hd__and3_2 _3461_ (
    .A(\g_bit[13].g_word[27].r_bit.Q ),
    .B(_0852_),
    .C(_0853_),
    .X(_1133_)
  );
  sky130_fd_sc_hd__a221o_2 _3462_ (
    .A1(\g_bit[13].g_word[6].r_bit.Q ),
    .A2(_0850_),
    .B1(_0851_),
    .B2(\g_bit[13].g_word[1].r_bit.Q ),
    .C1(_1133_),
    .X(_1134_)
  );
  sky130_fd_sc_hd__inv_2 _3463_ (
    .A(\g_bit[13].g_word[23].r_bit.Q ),
    .Y(_1135_)
  );
  sky130_fd_sc_hd__inv_2 _3464_ (
    .A(\g_bit[13].g_word[10].r_bit.Q ),
    .Y(_1136_)
  );
  sky130_fd_sc_hd__buf_1 _3465_ (
    .A(_0015_),
    .X(_1137_)
  );
  sky130_fd_sc_hd__or3_2 _3466_ (
    .A(_1136_),
    .B(_1137_),
    .C(_0700_),
    .X(_1138_)
  );
  sky130_fd_sc_hd__inv_2 _3467_ (
    .A(\g_bit[13].g_word[9].r_bit.Q ),
    .Y(_1139_)
  );
  sky130_fd_sc_hd__or3_2 _3468_ (
    .A(_1139_),
    .B(_0577_),
    .C(_0861_),
    .X(_1140_)
  );
  sky130_fd_sc_hd__inv_2 _3469_ (
    .A(\g_bit[13].g_word[8].r_bit.Q ),
    .Y(_1141_)
  );
  sky130_fd_sc_hd__or3_2 _3470_ (
    .A(_1141_),
    .B(_0705_),
    .C(_0864_),
    .X(_1142_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3471_ (
    .A1(_1135_),
    .A2(_0857_),
    .B1(_1138_),
    .C1(_1140_),
    .D1(_1142_),
    .Y(_1143_)
  );
  sky130_fd_sc_hd__inv_2 _3472_ (
    .A(\g_bit[13].g_word[22].r_bit.Q ),
    .Y(_1144_)
  );
  sky130_fd_sc_hd__inv_2 _3473_ (
    .A(\g_bit[13].g_word[16].r_bit.Q ),
    .Y(_1145_)
  );
  sky130_fd_sc_hd__or3_2 _3474_ (
    .A(_1145_),
    .B(_0584_),
    .C(_0870_),
    .X(_1146_)
  );
  sky130_fd_sc_hd__inv_2 _3475_ (
    .A(\g_bit[13].g_word[14].r_bit.Q ),
    .Y(_1147_)
  );
  sky130_fd_sc_hd__or3_2 _3476_ (
    .A(_1147_),
    .B(_0873_),
    .C(_0777_),
    .X(_1148_)
  );
  sky130_fd_sc_hd__inv_2 _3477_ (
    .A(\g_bit[13].g_word[18].r_bit.Q ),
    .Y(_1149_)
  );
  sky130_fd_sc_hd__or3_2 _3478_ (
    .A(_1149_),
    .B(_0780_),
    .C(_0876_),
    .X(_1150_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3479_ (
    .A1(_1144_),
    .A2(_0868_),
    .B1(_1146_),
    .C1(_1148_),
    .D1(_1150_),
    .Y(_1151_)
  );
  sky130_fd_sc_hd__or4_2 _3480_ (
    .A(_1132_),
    .B(_1134_),
    .C(_1143_),
    .D(_1151_),
    .X(_1152_)
  );
  sky130_fd_sc_hd__or4_2 _3481_ (
    .A(_1119_),
    .B(_1121_),
    .C(_1126_),
    .D(_1152_),
    .X(_1153_)
  );
  sky130_fd_sc_hd__buf_1 _3482_ (
    .A(_1153_),
    .X(\g_bit[13].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _3483_ (
    .A1(\g_bit[13].g_word[30].r_bit.Q ),
    .A2(_0883_),
    .A3(_0884_),
    .B1(_0885_),
    .B2(\g_bit[13].g_word[28].r_bit.Q ),
    .X(_1154_)
  );
  sky130_fd_sc_hd__a221o_2 _3484_ (
    .A1(\g_bit[13].g_word[4].r_bit.Q ),
    .A2(_0881_),
    .B1(_0882_),
    .B2(\g_bit[13].g_word[26].r_bit.Q ),
    .C1(_1154_),
    .X(_1155_)
  );
  sky130_fd_sc_hd__a22o_2 _3485_ (
    .A1(\g_bit[13].g_word[5].r_bit.Q ),
    .A2(_0890_),
    .B1(_0891_),
    .B2(\g_bit[13].g_word[2].r_bit.Q ),
    .X(_1156_)
  );
  sky130_fd_sc_hd__a221o_2 _3486_ (
    .A1(\g_bit[13].g_word[25].r_bit.Q ),
    .A2(_0888_),
    .B1(_0889_),
    .B2(\g_bit[13].g_word[31].r_bit.Q ),
    .C1(_1156_),
    .X(_1157_)
  );
  sky130_fd_sc_hd__a22o_2 _3487_ (
    .A1(\g_bit[13].g_word[13].r_bit.Q ),
    .A2(_0894_),
    .B1(_0895_),
    .B2(\g_bit[13].g_word[15].r_bit.Q ),
    .X(_1158_)
  );
  sky130_fd_sc_hd__a22o_2 _3488_ (
    .A1(\g_bit[13].g_word[20].r_bit.Q ),
    .A2(_0897_),
    .B1(_0898_),
    .B2(\g_bit[13].g_word[11].r_bit.Q ),
    .X(_1159_)
  );
  sky130_fd_sc_hd__a22o_2 _3489_ (
    .A1(\g_bit[13].g_word[19].r_bit.Q ),
    .A2(_0900_),
    .B1(_0901_),
    .B2(\g_bit[13].g_word[21].r_bit.Q ),
    .X(_1160_)
  );
  sky130_fd_sc_hd__a22o_2 _3490_ (
    .A1(\g_bit[13].g_word[17].r_bit.Q ),
    .A2(_0903_),
    .B1(_0904_),
    .B2(\g_bit[13].g_word[12].r_bit.Q ),
    .X(_1161_)
  );
  sky130_fd_sc_hd__or4_2 _3491_ (
    .A(_1158_),
    .B(_1159_),
    .C(_1160_),
    .D(_1161_),
    .X(_1162_)
  );
  sky130_fd_sc_hd__nor3_2 _3492_ (
    .A(_1127_),
    .B(_0794_),
    .C(_0727_),
    .Y(_1163_)
  );
  sky130_fd_sc_hd__nor3_2 _3493_ (
    .A(_1129_),
    .B(_0909_),
    .C(_0796_),
    .Y(_1164_)
  );
  sky130_fd_sc_hd__and3_2 _3494_ (
    .A(\g_bit[13].g_word[24].r_bit.Q ),
    .B(_0983_),
    .C(_0798_),
    .X(_1165_)
  );
  sky130_fd_sc_hd__a2111o_2 _3495_ (
    .A1(\g_bit[13].g_word[29].r_bit.Q ),
    .A2(_0907_),
    .B1(_1163_),
    .C1(_1164_),
    .D1(_1165_),
    .X(_1166_)
  );
  sky130_fd_sc_hd__and3_2 _3496_ (
    .A(\g_bit[13].g_word[27].r_bit.Q ),
    .B(_0915_),
    .C(_0916_),
    .X(_1167_)
  );
  sky130_fd_sc_hd__a221o_2 _3497_ (
    .A1(\g_bit[13].g_word[6].r_bit.Q ),
    .A2(_0913_),
    .B1(_0914_),
    .B2(\g_bit[13].g_word[1].r_bit.Q ),
    .C1(_1167_),
    .X(_1168_)
  );
  sky130_fd_sc_hd__buf_1 _3498_ (
    .A(_0144_),
    .X(_1169_)
  );
  sky130_fd_sc_hd__or3_2 _3499_ (
    .A(_1136_),
    .B(_1169_),
    .C(_0734_),
    .X(_1170_)
  );
  sky130_fd_sc_hd__or3_2 _3500_ (
    .A(_1139_),
    .B(_0609_),
    .C(_0921_),
    .X(_1171_)
  );
  sky130_fd_sc_hd__or3_2 _3501_ (
    .A(_1141_),
    .B(_0737_),
    .C(_0923_),
    .X(_1172_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3502_ (
    .A1(_1135_),
    .A2(_0919_),
    .B1(_1170_),
    .C1(_1171_),
    .D1(_1172_),
    .Y(_1173_)
  );
  sky130_fd_sc_hd__or3_2 _3503_ (
    .A(_1145_),
    .B(_0927_),
    .C(_0673_),
    .X(_1174_)
  );
  sky130_fd_sc_hd__or3_2 _3504_ (
    .A(_1147_),
    .B(_0929_),
    .C(_0808_),
    .X(_1175_)
  );
  sky130_fd_sc_hd__or3_2 _3505_ (
    .A(_1149_),
    .B(_0810_),
    .C(_0931_),
    .X(_1176_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3506_ (
    .A1(_1144_),
    .A2(_0926_),
    .B1(_1174_),
    .C1(_1175_),
    .D1(_1176_),
    .Y(_1177_)
  );
  sky130_fd_sc_hd__or4_2 _3507_ (
    .A(_1166_),
    .B(_1168_),
    .C(_1173_),
    .D(_1177_),
    .X(_1178_)
  );
  sky130_fd_sc_hd__or4_2 _3508_ (
    .A(_1155_),
    .B(_1157_),
    .C(_1162_),
    .D(_1178_),
    .X(_1179_)
  );
  sky130_fd_sc_hd__buf_1 _3509_ (
    .A(_1179_),
    .X(\g_bit[13].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _3510_ (
    .A1(\g_bit[14].g_word[30].r_bit.Q ),
    .A2(_0817_),
    .A3(_0818_),
    .B1(_0819_),
    .B2(\g_bit[14].g_word[28].r_bit.Q ),
    .X(_1180_)
  );
  sky130_fd_sc_hd__a221o_2 _3511_ (
    .A1(\g_bit[14].g_word[4].r_bit.Q ),
    .A2(_0815_),
    .B1(_0816_),
    .B2(\g_bit[14].g_word[26].r_bit.Q ),
    .C1(_1180_),
    .X(_1181_)
  );
  sky130_fd_sc_hd__a22o_2 _3512_ (
    .A1(\g_bit[14].g_word[5].r_bit.Q ),
    .A2(_0824_),
    .B1(_0825_),
    .B2(\g_bit[14].g_word[2].r_bit.Q ),
    .X(_1182_)
  );
  sky130_fd_sc_hd__a221o_2 _3513_ (
    .A1(\g_bit[14].g_word[25].r_bit.Q ),
    .A2(_0822_),
    .B1(_0823_),
    .B2(\g_bit[14].g_word[31].r_bit.Q ),
    .C1(_1182_),
    .X(_1183_)
  );
  sky130_fd_sc_hd__a22o_2 _3514_ (
    .A1(\g_bit[14].g_word[13].r_bit.Q ),
    .A2(_0828_),
    .B1(_0829_),
    .B2(\g_bit[14].g_word[15].r_bit.Q ),
    .X(_1184_)
  );
  sky130_fd_sc_hd__a22o_2 _3515_ (
    .A1(\g_bit[14].g_word[11].r_bit.Q ),
    .A2(_0831_),
    .B1(_0832_),
    .B2(\g_bit[14].g_word[20].r_bit.Q ),
    .X(_1185_)
  );
  sky130_fd_sc_hd__a22o_2 _3516_ (
    .A1(\g_bit[14].g_word[19].r_bit.Q ),
    .A2(_0834_),
    .B1(_0835_),
    .B2(\g_bit[14].g_word[21].r_bit.Q ),
    .X(_1186_)
  );
  sky130_fd_sc_hd__a22o_2 _3517_ (
    .A1(\g_bit[14].g_word[17].r_bit.Q ),
    .A2(_0837_),
    .B1(_0838_),
    .B2(\g_bit[14].g_word[12].r_bit.Q ),
    .X(_1187_)
  );
  sky130_fd_sc_hd__or4_2 _3518_ (
    .A(_1184_),
    .B(_1185_),
    .C(_1186_),
    .D(_1187_),
    .X(_1188_)
  );
  sky130_fd_sc_hd__inv_2 _3519_ (
    .A(\g_bit[14].g_word[7].r_bit.Q ),
    .Y(_1189_)
  );
  sky130_fd_sc_hd__nor3_2 _3520_ (
    .A(_1189_),
    .B(_0690_),
    .C(_0756_),
    .Y(_1190_)
  );
  sky130_fd_sc_hd__inv_2 _3521_ (
    .A(\g_bit[14].g_word[3].r_bit.Q ),
    .Y(_1191_)
  );
  sky130_fd_sc_hd__nor3_2 _3522_ (
    .A(_1191_),
    .B(_0845_),
    .C(_0846_),
    .Y(_1192_)
  );
  sky130_fd_sc_hd__and3_2 _3523_ (
    .A(\g_bit[14].g_word[24].r_bit.Q ),
    .B(_0760_),
    .C(_0949_),
    .X(_1193_)
  );
  sky130_fd_sc_hd__a2111o_2 _3524_ (
    .A1(\g_bit[14].g_word[29].r_bit.Q ),
    .A2(_0841_),
    .B1(_1190_),
    .C1(_1192_),
    .D1(_1193_),
    .X(_1194_)
  );
  sky130_fd_sc_hd__and3_2 _3525_ (
    .A(\g_bit[14].g_word[27].r_bit.Q ),
    .B(_0852_),
    .C(_0853_),
    .X(_1195_)
  );
  sky130_fd_sc_hd__a221o_2 _3526_ (
    .A1(\g_bit[14].g_word[6].r_bit.Q ),
    .A2(_0850_),
    .B1(_0851_),
    .B2(\g_bit[14].g_word[1].r_bit.Q ),
    .C1(_1195_),
    .X(_1196_)
  );
  sky130_fd_sc_hd__inv_2 _3527_ (
    .A(\g_bit[14].g_word[23].r_bit.Q ),
    .Y(_1197_)
  );
  sky130_fd_sc_hd__inv_2 _3528_ (
    .A(\g_bit[14].g_word[10].r_bit.Q ),
    .Y(_1198_)
  );
  sky130_fd_sc_hd__or3_2 _3529_ (
    .A(_1198_),
    .B(_1137_),
    .C(_0700_),
    .X(_1199_)
  );
  sky130_fd_sc_hd__inv_2 _3530_ (
    .A(\g_bit[14].g_word[9].r_bit.Q ),
    .Y(_1200_)
  );
  sky130_fd_sc_hd__or3_2 _3531_ (
    .A(_1200_),
    .B(_0577_),
    .C(_0861_),
    .X(_1201_)
  );
  sky130_fd_sc_hd__inv_2 _3532_ (
    .A(\g_bit[14].g_word[8].r_bit.Q ),
    .Y(_1202_)
  );
  sky130_fd_sc_hd__or3_2 _3533_ (
    .A(_1202_),
    .B(_0705_),
    .C(_0864_),
    .X(_1203_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3534_ (
    .A1(_1197_),
    .A2(_0857_),
    .B1(_1199_),
    .C1(_1201_),
    .D1(_1203_),
    .Y(_1204_)
  );
  sky130_fd_sc_hd__inv_2 _3535_ (
    .A(\g_bit[14].g_word[22].r_bit.Q ),
    .Y(_1205_)
  );
  sky130_fd_sc_hd__inv_2 _3536_ (
    .A(\g_bit[14].g_word[16].r_bit.Q ),
    .Y(_1206_)
  );
  sky130_fd_sc_hd__or3_2 _3537_ (
    .A(_1206_),
    .B(_0584_),
    .C(_0870_),
    .X(_1207_)
  );
  sky130_fd_sc_hd__inv_2 _3538_ (
    .A(\g_bit[14].g_word[14].r_bit.Q ),
    .Y(_1208_)
  );
  sky130_fd_sc_hd__or3_2 _3539_ (
    .A(_1208_),
    .B(_0873_),
    .C(_0777_),
    .X(_1209_)
  );
  sky130_fd_sc_hd__inv_2 _3540_ (
    .A(\g_bit[14].g_word[18].r_bit.Q ),
    .Y(_1210_)
  );
  sky130_fd_sc_hd__or3_2 _3541_ (
    .A(_1210_),
    .B(_0780_),
    .C(_0876_),
    .X(_1211_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3542_ (
    .A1(_1205_),
    .A2(_0868_),
    .B1(_1207_),
    .C1(_1209_),
    .D1(_1211_),
    .Y(_1212_)
  );
  sky130_fd_sc_hd__or4_2 _3543_ (
    .A(_1194_),
    .B(_1196_),
    .C(_1204_),
    .D(_1212_),
    .X(_1213_)
  );
  sky130_fd_sc_hd__or4_2 _3544_ (
    .A(_1181_),
    .B(_1183_),
    .C(_1188_),
    .D(_1213_),
    .X(_1214_)
  );
  sky130_fd_sc_hd__buf_1 _3545_ (
    .A(_1214_),
    .X(\g_bit[14].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _3546_ (
    .A1(\g_bit[14].g_word[30].r_bit.Q ),
    .A2(_0883_),
    .A3(_0884_),
    .B1(_0885_),
    .B2(\g_bit[14].g_word[28].r_bit.Q ),
    .X(_1215_)
  );
  sky130_fd_sc_hd__a221o_2 _3547_ (
    .A1(\g_bit[14].g_word[4].r_bit.Q ),
    .A2(_0881_),
    .B1(_0882_),
    .B2(\g_bit[14].g_word[26].r_bit.Q ),
    .C1(_1215_),
    .X(_1216_)
  );
  sky130_fd_sc_hd__a22o_2 _3548_ (
    .A1(\g_bit[14].g_word[5].r_bit.Q ),
    .A2(_0890_),
    .B1(_0891_),
    .B2(\g_bit[14].g_word[2].r_bit.Q ),
    .X(_1217_)
  );
  sky130_fd_sc_hd__a221o_2 _3549_ (
    .A1(\g_bit[14].g_word[25].r_bit.Q ),
    .A2(_0888_),
    .B1(_0889_),
    .B2(\g_bit[14].g_word[31].r_bit.Q ),
    .C1(_1217_),
    .X(_1218_)
  );
  sky130_fd_sc_hd__a22o_2 _3550_ (
    .A1(\g_bit[14].g_word[13].r_bit.Q ),
    .A2(_0894_),
    .B1(_0895_),
    .B2(\g_bit[14].g_word[15].r_bit.Q ),
    .X(_1219_)
  );
  sky130_fd_sc_hd__a22o_2 _3551_ (
    .A1(\g_bit[14].g_word[20].r_bit.Q ),
    .A2(_0897_),
    .B1(_0898_),
    .B2(\g_bit[14].g_word[11].r_bit.Q ),
    .X(_1220_)
  );
  sky130_fd_sc_hd__a22o_2 _3552_ (
    .A1(\g_bit[14].g_word[19].r_bit.Q ),
    .A2(_0900_),
    .B1(_0901_),
    .B2(\g_bit[14].g_word[21].r_bit.Q ),
    .X(_1221_)
  );
  sky130_fd_sc_hd__a22o_2 _3553_ (
    .A1(\g_bit[14].g_word[17].r_bit.Q ),
    .A2(_0903_),
    .B1(_0904_),
    .B2(\g_bit[14].g_word[12].r_bit.Q ),
    .X(_1222_)
  );
  sky130_fd_sc_hd__or4_2 _3554_ (
    .A(_1219_),
    .B(_1220_),
    .C(_1221_),
    .D(_1222_),
    .X(_1223_)
  );
  sky130_fd_sc_hd__nor3_2 _3555_ (
    .A(_1189_),
    .B(_0794_),
    .C(_0727_),
    .Y(_1224_)
  );
  sky130_fd_sc_hd__nor3_2 _3556_ (
    .A(_1191_),
    .B(_0909_),
    .C(_0796_),
    .Y(_1225_)
  );
  sky130_fd_sc_hd__and3_2 _3557_ (
    .A(\g_bit[14].g_word[24].r_bit.Q ),
    .B(_0983_),
    .C(_0798_),
    .X(_1226_)
  );
  sky130_fd_sc_hd__a2111o_2 _3558_ (
    .A1(\g_bit[14].g_word[29].r_bit.Q ),
    .A2(_0907_),
    .B1(_1224_),
    .C1(_1225_),
    .D1(_1226_),
    .X(_1227_)
  );
  sky130_fd_sc_hd__and3_2 _3559_ (
    .A(\g_bit[14].g_word[27].r_bit.Q ),
    .B(_0915_),
    .C(_0916_),
    .X(_1228_)
  );
  sky130_fd_sc_hd__a221o_2 _3560_ (
    .A1(\g_bit[14].g_word[6].r_bit.Q ),
    .A2(_0913_),
    .B1(_0914_),
    .B2(\g_bit[14].g_word[1].r_bit.Q ),
    .C1(_1228_),
    .X(_1229_)
  );
  sky130_fd_sc_hd__or3_2 _3561_ (
    .A(_1198_),
    .B(_1169_),
    .C(_0734_),
    .X(_1230_)
  );
  sky130_fd_sc_hd__or3_2 _3562_ (
    .A(_1200_),
    .B(_0609_),
    .C(_0921_),
    .X(_1231_)
  );
  sky130_fd_sc_hd__or3_2 _3563_ (
    .A(_1202_),
    .B(_0737_),
    .C(_0923_),
    .X(_1232_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3564_ (
    .A1(_1197_),
    .A2(_0919_),
    .B1(_1230_),
    .C1(_1231_),
    .D1(_1232_),
    .Y(_1233_)
  );
  sky130_fd_sc_hd__or3_2 _3565_ (
    .A(_1206_),
    .B(_0927_),
    .C(_0673_),
    .X(_1234_)
  );
  sky130_fd_sc_hd__or3_2 _3566_ (
    .A(_1208_),
    .B(_0929_),
    .C(_0808_),
    .X(_1235_)
  );
  sky130_fd_sc_hd__or3_2 _3567_ (
    .A(_1210_),
    .B(_0810_),
    .C(_0931_),
    .X(_1236_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3568_ (
    .A1(_1205_),
    .A2(_0926_),
    .B1(_1234_),
    .C1(_1235_),
    .D1(_1236_),
    .Y(_1237_)
  );
  sky130_fd_sc_hd__or4_2 _3569_ (
    .A(_1227_),
    .B(_1229_),
    .C(_1233_),
    .D(_1237_),
    .X(_1238_)
  );
  sky130_fd_sc_hd__or4_2 _3570_ (
    .A(_1216_),
    .B(_1218_),
    .C(_1223_),
    .D(_1238_),
    .X(_1239_)
  );
  sky130_fd_sc_hd__buf_1 _3571_ (
    .A(_1239_),
    .X(\g_bit[14].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _3572_ (
    .A1(\g_bit[15].g_word[30].r_bit.Q ),
    .A2(_0817_),
    .A3(_0818_),
    .B1(_0819_),
    .B2(\g_bit[15].g_word[28].r_bit.Q ),
    .X(_1240_)
  );
  sky130_fd_sc_hd__a221o_2 _3573_ (
    .A1(\g_bit[15].g_word[4].r_bit.Q ),
    .A2(_0815_),
    .B1(_0816_),
    .B2(\g_bit[15].g_word[26].r_bit.Q ),
    .C1(_1240_),
    .X(_1241_)
  );
  sky130_fd_sc_hd__a22o_2 _3574_ (
    .A1(\g_bit[15].g_word[5].r_bit.Q ),
    .A2(_0824_),
    .B1(_0825_),
    .B2(\g_bit[15].g_word[2].r_bit.Q ),
    .X(_1242_)
  );
  sky130_fd_sc_hd__a221o_2 _3575_ (
    .A1(\g_bit[15].g_word[25].r_bit.Q ),
    .A2(_0822_),
    .B1(_0823_),
    .B2(\g_bit[15].g_word[31].r_bit.Q ),
    .C1(_1242_),
    .X(_1243_)
  );
  sky130_fd_sc_hd__a22o_2 _3576_ (
    .A1(\g_bit[15].g_word[13].r_bit.Q ),
    .A2(_0828_),
    .B1(_0829_),
    .B2(\g_bit[15].g_word[15].r_bit.Q ),
    .X(_1244_)
  );
  sky130_fd_sc_hd__a22o_2 _3577_ (
    .A1(\g_bit[15].g_word[11].r_bit.Q ),
    .A2(_0831_),
    .B1(_0832_),
    .B2(\g_bit[15].g_word[20].r_bit.Q ),
    .X(_1245_)
  );
  sky130_fd_sc_hd__a22o_2 _3578_ (
    .A1(\g_bit[15].g_word[19].r_bit.Q ),
    .A2(_0834_),
    .B1(_0835_),
    .B2(\g_bit[15].g_word[21].r_bit.Q ),
    .X(_1246_)
  );
  sky130_fd_sc_hd__a22o_2 _3579_ (
    .A1(\g_bit[15].g_word[17].r_bit.Q ),
    .A2(_0837_),
    .B1(_0838_),
    .B2(\g_bit[15].g_word[12].r_bit.Q ),
    .X(_1247_)
  );
  sky130_fd_sc_hd__or4_2 _3580_ (
    .A(_1244_),
    .B(_1245_),
    .C(_1246_),
    .D(_1247_),
    .X(_1248_)
  );
  sky130_fd_sc_hd__inv_2 _3581_ (
    .A(\g_bit[15].g_word[7].r_bit.Q ),
    .Y(_1249_)
  );
  sky130_fd_sc_hd__nor3_2 _3582_ (
    .A(_1249_),
    .B(_0690_),
    .C(_0756_),
    .Y(_1250_)
  );
  sky130_fd_sc_hd__inv_2 _3583_ (
    .A(\g_bit[15].g_word[3].r_bit.Q ),
    .Y(_1251_)
  );
  sky130_fd_sc_hd__nor3_2 _3584_ (
    .A(_1251_),
    .B(_0845_),
    .C(_0846_),
    .Y(_1252_)
  );
  sky130_fd_sc_hd__and3_2 _3585_ (
    .A(\g_bit[15].g_word[24].r_bit.Q ),
    .B(_0760_),
    .C(_0949_),
    .X(_1253_)
  );
  sky130_fd_sc_hd__a2111o_2 _3586_ (
    .A1(\g_bit[15].g_word[29].r_bit.Q ),
    .A2(_0841_),
    .B1(_1250_),
    .C1(_1252_),
    .D1(_1253_),
    .X(_1254_)
  );
  sky130_fd_sc_hd__and3_2 _3587_ (
    .A(\g_bit[15].g_word[27].r_bit.Q ),
    .B(_0852_),
    .C(_0853_),
    .X(_1255_)
  );
  sky130_fd_sc_hd__a221o_2 _3588_ (
    .A1(\g_bit[15].g_word[6].r_bit.Q ),
    .A2(_0850_),
    .B1(_0851_),
    .B2(\g_bit[15].g_word[1].r_bit.Q ),
    .C1(_1255_),
    .X(_1256_)
  );
  sky130_fd_sc_hd__inv_2 _3589_ (
    .A(\g_bit[15].g_word[23].r_bit.Q ),
    .Y(_1257_)
  );
  sky130_fd_sc_hd__inv_2 _3590_ (
    .A(\g_bit[15].g_word[10].r_bit.Q ),
    .Y(_1258_)
  );
  sky130_fd_sc_hd__or3_2 _3591_ (
    .A(_1258_),
    .B(_1137_),
    .C(_0700_),
    .X(_1259_)
  );
  sky130_fd_sc_hd__inv_2 _3592_ (
    .A(\g_bit[15].g_word[9].r_bit.Q ),
    .Y(_1260_)
  );
  sky130_fd_sc_hd__buf_1 _3593_ (
    .A(_0015_),
    .X(_1261_)
  );
  sky130_fd_sc_hd__or3_2 _3594_ (
    .A(_1260_),
    .B(_1261_),
    .C(_0861_),
    .X(_1262_)
  );
  sky130_fd_sc_hd__inv_2 _3595_ (
    .A(\g_bit[15].g_word[8].r_bit.Q ),
    .Y(_1263_)
  );
  sky130_fd_sc_hd__or3_2 _3596_ (
    .A(_1263_),
    .B(_0705_),
    .C(_0864_),
    .X(_1264_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3597_ (
    .A1(_1257_),
    .A2(_0857_),
    .B1(_1259_),
    .C1(_1262_),
    .D1(_1264_),
    .Y(_1265_)
  );
  sky130_fd_sc_hd__inv_2 _3598_ (
    .A(\g_bit[15].g_word[22].r_bit.Q ),
    .Y(_1266_)
  );
  sky130_fd_sc_hd__inv_2 _3599_ (
    .A(\g_bit[15].g_word[16].r_bit.Q ),
    .Y(_1267_)
  );
  sky130_fd_sc_hd__buf_1 _3600_ (
    .A(_0045_),
    .X(_1268_)
  );
  sky130_fd_sc_hd__or3_2 _3601_ (
    .A(_1267_),
    .B(_1268_),
    .C(_0870_),
    .X(_1269_)
  );
  sky130_fd_sc_hd__inv_2 _3602_ (
    .A(\g_bit[15].g_word[14].r_bit.Q ),
    .Y(_1270_)
  );
  sky130_fd_sc_hd__or3_2 _3603_ (
    .A(_1270_),
    .B(_0873_),
    .C(_0777_),
    .X(_1271_)
  );
  sky130_fd_sc_hd__inv_2 _3604_ (
    .A(\g_bit[15].g_word[18].r_bit.Q ),
    .Y(_1272_)
  );
  sky130_fd_sc_hd__or3_2 _3605_ (
    .A(_1272_),
    .B(_0780_),
    .C(_0876_),
    .X(_1273_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3606_ (
    .A1(_1266_),
    .A2(_0868_),
    .B1(_1269_),
    .C1(_1271_),
    .D1(_1273_),
    .Y(_1274_)
  );
  sky130_fd_sc_hd__or4_2 _3607_ (
    .A(_1254_),
    .B(_1256_),
    .C(_1265_),
    .D(_1274_),
    .X(_1275_)
  );
  sky130_fd_sc_hd__or4_2 _3608_ (
    .A(_1241_),
    .B(_1243_),
    .C(_1248_),
    .D(_1275_),
    .X(_1276_)
  );
  sky130_fd_sc_hd__buf_1 _3609_ (
    .A(_1276_),
    .X(\g_bit[15].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _3610_ (
    .A1(\g_bit[15].g_word[30].r_bit.Q ),
    .A2(_0883_),
    .A3(_0884_),
    .B1(_0885_),
    .B2(\g_bit[15].g_word[28].r_bit.Q ),
    .X(_1277_)
  );
  sky130_fd_sc_hd__a221o_2 _3611_ (
    .A1(\g_bit[15].g_word[4].r_bit.Q ),
    .A2(_0881_),
    .B1(_0882_),
    .B2(\g_bit[15].g_word[26].r_bit.Q ),
    .C1(_1277_),
    .X(_1278_)
  );
  sky130_fd_sc_hd__a22o_2 _3612_ (
    .A1(\g_bit[15].g_word[5].r_bit.Q ),
    .A2(_0890_),
    .B1(_0891_),
    .B2(\g_bit[15].g_word[2].r_bit.Q ),
    .X(_1279_)
  );
  sky130_fd_sc_hd__a221o_2 _3613_ (
    .A1(\g_bit[15].g_word[25].r_bit.Q ),
    .A2(_0888_),
    .B1(_0889_),
    .B2(\g_bit[15].g_word[31].r_bit.Q ),
    .C1(_1279_),
    .X(_1280_)
  );
  sky130_fd_sc_hd__a22o_2 _3614_ (
    .A1(\g_bit[15].g_word[13].r_bit.Q ),
    .A2(_0894_),
    .B1(_0895_),
    .B2(\g_bit[15].g_word[15].r_bit.Q ),
    .X(_1281_)
  );
  sky130_fd_sc_hd__a22o_2 _3615_ (
    .A1(\g_bit[15].g_word[20].r_bit.Q ),
    .A2(_0897_),
    .B1(_0898_),
    .B2(\g_bit[15].g_word[11].r_bit.Q ),
    .X(_1282_)
  );
  sky130_fd_sc_hd__a22o_2 _3616_ (
    .A1(\g_bit[15].g_word[19].r_bit.Q ),
    .A2(_0900_),
    .B1(_0901_),
    .B2(\g_bit[15].g_word[21].r_bit.Q ),
    .X(_1283_)
  );
  sky130_fd_sc_hd__a22o_2 _3617_ (
    .A1(\g_bit[15].g_word[17].r_bit.Q ),
    .A2(_0903_),
    .B1(_0904_),
    .B2(\g_bit[15].g_word[12].r_bit.Q ),
    .X(_1284_)
  );
  sky130_fd_sc_hd__or4_2 _3618_ (
    .A(_1281_),
    .B(_1282_),
    .C(_1283_),
    .D(_1284_),
    .X(_1285_)
  );
  sky130_fd_sc_hd__nor3_2 _3619_ (
    .A(_1249_),
    .B(_0794_),
    .C(_0727_),
    .Y(_1286_)
  );
  sky130_fd_sc_hd__nor3_2 _3620_ (
    .A(_1251_),
    .B(_0909_),
    .C(_0796_),
    .Y(_1287_)
  );
  sky130_fd_sc_hd__and3_2 _3621_ (
    .A(\g_bit[15].g_word[24].r_bit.Q ),
    .B(_0983_),
    .C(_0798_),
    .X(_1288_)
  );
  sky130_fd_sc_hd__a2111o_2 _3622_ (
    .A1(\g_bit[15].g_word[29].r_bit.Q ),
    .A2(_0907_),
    .B1(_1286_),
    .C1(_1287_),
    .D1(_1288_),
    .X(_1289_)
  );
  sky130_fd_sc_hd__and3_2 _3623_ (
    .A(\g_bit[15].g_word[27].r_bit.Q ),
    .B(_0915_),
    .C(_0916_),
    .X(_1290_)
  );
  sky130_fd_sc_hd__a221o_2 _3624_ (
    .A1(\g_bit[15].g_word[6].r_bit.Q ),
    .A2(_0913_),
    .B1(_0914_),
    .B2(\g_bit[15].g_word[1].r_bit.Q ),
    .C1(_1290_),
    .X(_1291_)
  );
  sky130_fd_sc_hd__or3_2 _3625_ (
    .A(_1258_),
    .B(_1169_),
    .C(_0734_),
    .X(_1292_)
  );
  sky130_fd_sc_hd__buf_1 _3626_ (
    .A(_0144_),
    .X(_1293_)
  );
  sky130_fd_sc_hd__or3_2 _3627_ (
    .A(_1260_),
    .B(_1293_),
    .C(_0921_),
    .X(_1294_)
  );
  sky130_fd_sc_hd__or3_2 _3628_ (
    .A(_1263_),
    .B(_0737_),
    .C(_0923_),
    .X(_1295_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3629_ (
    .A1(_1257_),
    .A2(_0919_),
    .B1(_1292_),
    .C1(_1294_),
    .D1(_1295_),
    .Y(_1296_)
  );
  sky130_fd_sc_hd__or3_2 _3630_ (
    .A(_1267_),
    .B(_0927_),
    .C(_0673_),
    .X(_1297_)
  );
  sky130_fd_sc_hd__or3_2 _3631_ (
    .A(_1270_),
    .B(_0929_),
    .C(_0808_),
    .X(_1298_)
  );
  sky130_fd_sc_hd__or3_2 _3632_ (
    .A(_1272_),
    .B(_0810_),
    .C(_0931_),
    .X(_1299_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3633_ (
    .A1(_1266_),
    .A2(_0926_),
    .B1(_1297_),
    .C1(_1298_),
    .D1(_1299_),
    .Y(_1300_)
  );
  sky130_fd_sc_hd__or4_2 _3634_ (
    .A(_1289_),
    .B(_1291_),
    .C(_1296_),
    .D(_1300_),
    .X(_1301_)
  );
  sky130_fd_sc_hd__or4_2 _3635_ (
    .A(_1278_),
    .B(_1280_),
    .C(_1285_),
    .D(_1301_),
    .X(_1302_)
  );
  sky130_fd_sc_hd__buf_1 _3636_ (
    .A(_1302_),
    .X(\g_bit[15].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _3637_ (
    .A1(\g_bit[16].g_word[30].r_bit.Q ),
    .A2(_0817_),
    .A3(_0818_),
    .B1(_0819_),
    .B2(\g_bit[16].g_word[28].r_bit.Q ),
    .X(_1303_)
  );
  sky130_fd_sc_hd__a221o_2 _3638_ (
    .A1(\g_bit[16].g_word[4].r_bit.Q ),
    .A2(_0815_),
    .B1(_0816_),
    .B2(\g_bit[16].g_word[26].r_bit.Q ),
    .C1(_1303_),
    .X(_1304_)
  );
  sky130_fd_sc_hd__a22o_2 _3639_ (
    .A1(\g_bit[16].g_word[5].r_bit.Q ),
    .A2(_0824_),
    .B1(_0825_),
    .B2(\g_bit[16].g_word[2].r_bit.Q ),
    .X(_1305_)
  );
  sky130_fd_sc_hd__a221o_2 _3640_ (
    .A1(\g_bit[16].g_word[25].r_bit.Q ),
    .A2(_0822_),
    .B1(_0823_),
    .B2(\g_bit[16].g_word[31].r_bit.Q ),
    .C1(_1305_),
    .X(_1306_)
  );
  sky130_fd_sc_hd__a22o_2 _3641_ (
    .A1(\g_bit[16].g_word[13].r_bit.Q ),
    .A2(_0828_),
    .B1(_0829_),
    .B2(\g_bit[16].g_word[15].r_bit.Q ),
    .X(_1307_)
  );
  sky130_fd_sc_hd__a22o_2 _3642_ (
    .A1(\g_bit[16].g_word[11].r_bit.Q ),
    .A2(_0831_),
    .B1(_0832_),
    .B2(\g_bit[16].g_word[20].r_bit.Q ),
    .X(_1308_)
  );
  sky130_fd_sc_hd__a22o_2 _3643_ (
    .A1(\g_bit[16].g_word[19].r_bit.Q ),
    .A2(_0834_),
    .B1(_0835_),
    .B2(\g_bit[16].g_word[21].r_bit.Q ),
    .X(_1309_)
  );
  sky130_fd_sc_hd__a22o_2 _3644_ (
    .A1(\g_bit[16].g_word[17].r_bit.Q ),
    .A2(_0837_),
    .B1(_0838_),
    .B2(\g_bit[16].g_word[12].r_bit.Q ),
    .X(_1310_)
  );
  sky130_fd_sc_hd__or4_2 _3645_ (
    .A(_1307_),
    .B(_1308_),
    .C(_1309_),
    .D(_1310_),
    .X(_1311_)
  );
  sky130_fd_sc_hd__inv_2 _3646_ (
    .A(\g_bit[16].g_word[7].r_bit.Q ),
    .Y(_1312_)
  );
  sky130_fd_sc_hd__nor3_2 _3647_ (
    .A(_1312_),
    .B(_0690_),
    .C(_0756_),
    .Y(_1313_)
  );
  sky130_fd_sc_hd__inv_2 _3648_ (
    .A(\g_bit[16].g_word[3].r_bit.Q ),
    .Y(_1314_)
  );
  sky130_fd_sc_hd__nor3_2 _3649_ (
    .A(_1314_),
    .B(_0845_),
    .C(_0846_),
    .Y(_1315_)
  );
  sky130_fd_sc_hd__and3_2 _3650_ (
    .A(\g_bit[16].g_word[24].r_bit.Q ),
    .B(_0760_),
    .C(_0949_),
    .X(_1316_)
  );
  sky130_fd_sc_hd__a2111o_2 _3651_ (
    .A1(\g_bit[16].g_word[29].r_bit.Q ),
    .A2(_0841_),
    .B1(_1313_),
    .C1(_1315_),
    .D1(_1316_),
    .X(_1317_)
  );
  sky130_fd_sc_hd__and3_2 _3652_ (
    .A(\g_bit[16].g_word[27].r_bit.Q ),
    .B(_0852_),
    .C(_0853_),
    .X(_1318_)
  );
  sky130_fd_sc_hd__a221o_2 _3653_ (
    .A1(\g_bit[16].g_word[6].r_bit.Q ),
    .A2(_0850_),
    .B1(_0851_),
    .B2(\g_bit[16].g_word[1].r_bit.Q ),
    .C1(_1318_),
    .X(_1319_)
  );
  sky130_fd_sc_hd__inv_2 _3654_ (
    .A(\g_bit[16].g_word[23].r_bit.Q ),
    .Y(_1320_)
  );
  sky130_fd_sc_hd__inv_2 _3655_ (
    .A(\g_bit[16].g_word[10].r_bit.Q ),
    .Y(_1321_)
  );
  sky130_fd_sc_hd__or3_2 _3656_ (
    .A(_1321_),
    .B(_1137_),
    .C(_0700_),
    .X(_1322_)
  );
  sky130_fd_sc_hd__inv_2 _3657_ (
    .A(\g_bit[16].g_word[9].r_bit.Q ),
    .Y(_1323_)
  );
  sky130_fd_sc_hd__or3_2 _3658_ (
    .A(_1323_),
    .B(_1261_),
    .C(_0861_),
    .X(_1324_)
  );
  sky130_fd_sc_hd__inv_2 _3659_ (
    .A(\g_bit[16].g_word[8].r_bit.Q ),
    .Y(_1325_)
  );
  sky130_fd_sc_hd__or3_2 _3660_ (
    .A(_1325_),
    .B(_0705_),
    .C(_0864_),
    .X(_1326_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3661_ (
    .A1(_1320_),
    .A2(_0857_),
    .B1(_1322_),
    .C1(_1324_),
    .D1(_1326_),
    .Y(_1327_)
  );
  sky130_fd_sc_hd__inv_2 _3662_ (
    .A(\g_bit[16].g_word[22].r_bit.Q ),
    .Y(_1328_)
  );
  sky130_fd_sc_hd__inv_2 _3663_ (
    .A(\g_bit[16].g_word[16].r_bit.Q ),
    .Y(_1329_)
  );
  sky130_fd_sc_hd__or3_2 _3664_ (
    .A(_1329_),
    .B(_1268_),
    .C(_0870_),
    .X(_1330_)
  );
  sky130_fd_sc_hd__inv_2 _3665_ (
    .A(\g_bit[16].g_word[14].r_bit.Q ),
    .Y(_1331_)
  );
  sky130_fd_sc_hd__or3_2 _3666_ (
    .A(_1331_),
    .B(_0873_),
    .C(_0777_),
    .X(_1332_)
  );
  sky130_fd_sc_hd__inv_2 _3667_ (
    .A(\g_bit[16].g_word[18].r_bit.Q ),
    .Y(_1333_)
  );
  sky130_fd_sc_hd__or3_2 _3668_ (
    .A(_1333_),
    .B(_0780_),
    .C(_0876_),
    .X(_1334_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3669_ (
    .A1(_1328_),
    .A2(_0868_),
    .B1(_1330_),
    .C1(_1332_),
    .D1(_1334_),
    .Y(_1335_)
  );
  sky130_fd_sc_hd__or4_2 _3670_ (
    .A(_1317_),
    .B(_1319_),
    .C(_1327_),
    .D(_1335_),
    .X(_1336_)
  );
  sky130_fd_sc_hd__or4_2 _3671_ (
    .A(_1304_),
    .B(_1306_),
    .C(_1311_),
    .D(_1336_),
    .X(_1337_)
  );
  sky130_fd_sc_hd__buf_1 _3672_ (
    .A(_1337_),
    .X(\g_bit[16].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _3673_ (
    .A1(\g_bit[16].g_word[30].r_bit.Q ),
    .A2(_0883_),
    .A3(_0884_),
    .B1(_0885_),
    .B2(\g_bit[16].g_word[28].r_bit.Q ),
    .X(_1338_)
  );
  sky130_fd_sc_hd__a221o_2 _3674_ (
    .A1(\g_bit[16].g_word[4].r_bit.Q ),
    .A2(_0881_),
    .B1(_0882_),
    .B2(\g_bit[16].g_word[26].r_bit.Q ),
    .C1(_1338_),
    .X(_1339_)
  );
  sky130_fd_sc_hd__a22o_2 _3675_ (
    .A1(\g_bit[16].g_word[5].r_bit.Q ),
    .A2(_0890_),
    .B1(_0891_),
    .B2(\g_bit[16].g_word[2].r_bit.Q ),
    .X(_1340_)
  );
  sky130_fd_sc_hd__a221o_2 _3676_ (
    .A1(\g_bit[16].g_word[25].r_bit.Q ),
    .A2(_0888_),
    .B1(_0889_),
    .B2(\g_bit[16].g_word[31].r_bit.Q ),
    .C1(_1340_),
    .X(_1341_)
  );
  sky130_fd_sc_hd__a22o_2 _3677_ (
    .A1(\g_bit[16].g_word[13].r_bit.Q ),
    .A2(_0894_),
    .B1(_0895_),
    .B2(\g_bit[16].g_word[15].r_bit.Q ),
    .X(_1342_)
  );
  sky130_fd_sc_hd__a22o_2 _3678_ (
    .A1(\g_bit[16].g_word[20].r_bit.Q ),
    .A2(_0897_),
    .B1(_0898_),
    .B2(\g_bit[16].g_word[11].r_bit.Q ),
    .X(_1343_)
  );
  sky130_fd_sc_hd__a22o_2 _3679_ (
    .A1(\g_bit[16].g_word[19].r_bit.Q ),
    .A2(_0900_),
    .B1(_0901_),
    .B2(\g_bit[16].g_word[21].r_bit.Q ),
    .X(_1344_)
  );
  sky130_fd_sc_hd__a22o_2 _3680_ (
    .A1(\g_bit[16].g_word[17].r_bit.Q ),
    .A2(_0903_),
    .B1(_0904_),
    .B2(\g_bit[16].g_word[12].r_bit.Q ),
    .X(_1345_)
  );
  sky130_fd_sc_hd__or4_2 _3681_ (
    .A(_1342_),
    .B(_1343_),
    .C(_1344_),
    .D(_1345_),
    .X(_1346_)
  );
  sky130_fd_sc_hd__nor3_2 _3682_ (
    .A(_1312_),
    .B(_0794_),
    .C(_0727_),
    .Y(_1347_)
  );
  sky130_fd_sc_hd__nor3_2 _3683_ (
    .A(_1314_),
    .B(_0909_),
    .C(_0796_),
    .Y(_1348_)
  );
  sky130_fd_sc_hd__and3_2 _3684_ (
    .A(\g_bit[16].g_word[24].r_bit.Q ),
    .B(_0983_),
    .C(_0798_),
    .X(_1349_)
  );
  sky130_fd_sc_hd__a2111o_2 _3685_ (
    .A1(\g_bit[16].g_word[29].r_bit.Q ),
    .A2(_0907_),
    .B1(_1347_),
    .C1(_1348_),
    .D1(_1349_),
    .X(_1350_)
  );
  sky130_fd_sc_hd__and3_2 _3686_ (
    .A(\g_bit[16].g_word[27].r_bit.Q ),
    .B(_0915_),
    .C(_0916_),
    .X(_1351_)
  );
  sky130_fd_sc_hd__a221o_2 _3687_ (
    .A1(\g_bit[16].g_word[6].r_bit.Q ),
    .A2(_0913_),
    .B1(_0914_),
    .B2(\g_bit[16].g_word[1].r_bit.Q ),
    .C1(_1351_),
    .X(_1352_)
  );
  sky130_fd_sc_hd__or3_2 _3688_ (
    .A(_1321_),
    .B(_1169_),
    .C(_0734_),
    .X(_1353_)
  );
  sky130_fd_sc_hd__or3_2 _3689_ (
    .A(_1323_),
    .B(_1293_),
    .C(_0921_),
    .X(_1354_)
  );
  sky130_fd_sc_hd__or3_2 _3690_ (
    .A(_1325_),
    .B(_0737_),
    .C(_0923_),
    .X(_1355_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3691_ (
    .A1(_1320_),
    .A2(_0919_),
    .B1(_1353_),
    .C1(_1354_),
    .D1(_1355_),
    .Y(_1356_)
  );
  sky130_fd_sc_hd__buf_1 _3692_ (
    .A(_0174_),
    .X(_1357_)
  );
  sky130_fd_sc_hd__or3_2 _3693_ (
    .A(_1329_),
    .B(_0927_),
    .C(_1357_),
    .X(_1358_)
  );
  sky130_fd_sc_hd__or3_2 _3694_ (
    .A(_1331_),
    .B(_0929_),
    .C(_0808_),
    .X(_1359_)
  );
  sky130_fd_sc_hd__or3_2 _3695_ (
    .A(_1333_),
    .B(_0810_),
    .C(_0931_),
    .X(_1360_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3696_ (
    .A1(_1328_),
    .A2(_0926_),
    .B1(_1358_),
    .C1(_1359_),
    .D1(_1360_),
    .Y(_1361_)
  );
  sky130_fd_sc_hd__or4_2 _3697_ (
    .A(_1350_),
    .B(_1352_),
    .C(_1356_),
    .D(_1361_),
    .X(_1362_)
  );
  sky130_fd_sc_hd__or4_2 _3698_ (
    .A(_1339_),
    .B(_1341_),
    .C(_1346_),
    .D(_1362_),
    .X(_1363_)
  );
  sky130_fd_sc_hd__buf_1 _3699_ (
    .A(_1363_),
    .X(\g_bit[16].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _3700_ (
    .A1(\g_bit[17].g_word[30].r_bit.Q ),
    .A2(_0817_),
    .A3(_0818_),
    .B1(_0819_),
    .B2(\g_bit[17].g_word[28].r_bit.Q ),
    .X(_1364_)
  );
  sky130_fd_sc_hd__a221o_2 _3701_ (
    .A1(\g_bit[17].g_word[4].r_bit.Q ),
    .A2(_0815_),
    .B1(_0816_),
    .B2(\g_bit[17].g_word[26].r_bit.Q ),
    .C1(_1364_),
    .X(_1365_)
  );
  sky130_fd_sc_hd__a22o_2 _3702_ (
    .A1(\g_bit[17].g_word[5].r_bit.Q ),
    .A2(_0824_),
    .B1(_0825_),
    .B2(\g_bit[17].g_word[2].r_bit.Q ),
    .X(_1366_)
  );
  sky130_fd_sc_hd__a221o_2 _3703_ (
    .A1(\g_bit[17].g_word[25].r_bit.Q ),
    .A2(_0822_),
    .B1(_0823_),
    .B2(\g_bit[17].g_word[31].r_bit.Q ),
    .C1(_1366_),
    .X(_1367_)
  );
  sky130_fd_sc_hd__a22o_2 _3704_ (
    .A1(\g_bit[17].g_word[13].r_bit.Q ),
    .A2(_0828_),
    .B1(_0829_),
    .B2(\g_bit[17].g_word[15].r_bit.Q ),
    .X(_1368_)
  );
  sky130_fd_sc_hd__a22o_2 _3705_ (
    .A1(\g_bit[17].g_word[11].r_bit.Q ),
    .A2(_0831_),
    .B1(_0832_),
    .B2(\g_bit[17].g_word[20].r_bit.Q ),
    .X(_1369_)
  );
  sky130_fd_sc_hd__a22o_2 _3706_ (
    .A1(\g_bit[17].g_word[19].r_bit.Q ),
    .A2(_0834_),
    .B1(_0835_),
    .B2(\g_bit[17].g_word[21].r_bit.Q ),
    .X(_1370_)
  );
  sky130_fd_sc_hd__a22o_2 _3707_ (
    .A1(\g_bit[17].g_word[17].r_bit.Q ),
    .A2(_0837_),
    .B1(_0838_),
    .B2(\g_bit[17].g_word[12].r_bit.Q ),
    .X(_1371_)
  );
  sky130_fd_sc_hd__or4_2 _3708_ (
    .A(_1368_),
    .B(_1369_),
    .C(_1370_),
    .D(_1371_),
    .X(_1372_)
  );
  sky130_fd_sc_hd__inv_2 _3709_ (
    .A(\g_bit[17].g_word[7].r_bit.Q ),
    .Y(_1373_)
  );
  sky130_fd_sc_hd__buf_1 _3710_ (
    .A(_0081_),
    .X(_1374_)
  );
  sky130_fd_sc_hd__nor3_2 _3711_ (
    .A(_1373_),
    .B(_1374_),
    .C(_0756_),
    .Y(_1375_)
  );
  sky130_fd_sc_hd__inv_2 _3712_ (
    .A(\g_bit[17].g_word[3].r_bit.Q ),
    .Y(_1376_)
  );
  sky130_fd_sc_hd__nor3_2 _3713_ (
    .A(_1376_),
    .B(_0845_),
    .C(_0846_),
    .Y(_1377_)
  );
  sky130_fd_sc_hd__and3_2 _3714_ (
    .A(\g_bit[17].g_word[24].r_bit.Q ),
    .B(_0760_),
    .C(_0949_),
    .X(_1378_)
  );
  sky130_fd_sc_hd__a2111o_2 _3715_ (
    .A1(\g_bit[17].g_word[29].r_bit.Q ),
    .A2(_0841_),
    .B1(_1375_),
    .C1(_1377_),
    .D1(_1378_),
    .X(_1379_)
  );
  sky130_fd_sc_hd__and3_2 _3716_ (
    .A(\g_bit[17].g_word[27].r_bit.Q ),
    .B(_0852_),
    .C(_0853_),
    .X(_1380_)
  );
  sky130_fd_sc_hd__a221o_2 _3717_ (
    .A1(\g_bit[17].g_word[6].r_bit.Q ),
    .A2(_0850_),
    .B1(_0851_),
    .B2(\g_bit[17].g_word[1].r_bit.Q ),
    .C1(_1380_),
    .X(_1381_)
  );
  sky130_fd_sc_hd__inv_2 _3718_ (
    .A(\g_bit[17].g_word[23].r_bit.Q ),
    .Y(_1382_)
  );
  sky130_fd_sc_hd__inv_2 _3719_ (
    .A(\g_bit[17].g_word[10].r_bit.Q ),
    .Y(_1383_)
  );
  sky130_fd_sc_hd__buf_1 _3720_ (
    .A(_0048_),
    .X(_1384_)
  );
  sky130_fd_sc_hd__or3_2 _3721_ (
    .A(_1383_),
    .B(_1137_),
    .C(_1384_),
    .X(_1385_)
  );
  sky130_fd_sc_hd__inv_2 _3722_ (
    .A(\g_bit[17].g_word[9].r_bit.Q ),
    .Y(_1386_)
  );
  sky130_fd_sc_hd__or3_2 _3723_ (
    .A(_1386_),
    .B(_1261_),
    .C(_0861_),
    .X(_1387_)
  );
  sky130_fd_sc_hd__inv_2 _3724_ (
    .A(\g_bit[17].g_word[8].r_bit.Q ),
    .Y(_1388_)
  );
  sky130_fd_sc_hd__buf_1 _3725_ (
    .A(_0015_),
    .X(_1389_)
  );
  sky130_fd_sc_hd__or3_2 _3726_ (
    .A(_1388_),
    .B(_1389_),
    .C(_0864_),
    .X(_1390_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3727_ (
    .A1(_1382_),
    .A2(_0857_),
    .B1(_1385_),
    .C1(_1387_),
    .D1(_1390_),
    .Y(_1391_)
  );
  sky130_fd_sc_hd__inv_2 _3728_ (
    .A(\g_bit[17].g_word[22].r_bit.Q ),
    .Y(_1392_)
  );
  sky130_fd_sc_hd__inv_2 _3729_ (
    .A(\g_bit[17].g_word[16].r_bit.Q ),
    .Y(_1393_)
  );
  sky130_fd_sc_hd__or3_2 _3730_ (
    .A(_1393_),
    .B(_1268_),
    .C(_0870_),
    .X(_1394_)
  );
  sky130_fd_sc_hd__inv_2 _3731_ (
    .A(\g_bit[17].g_word[14].r_bit.Q ),
    .Y(_1395_)
  );
  sky130_fd_sc_hd__or3_2 _3732_ (
    .A(_1395_),
    .B(_0873_),
    .C(_0777_),
    .X(_1396_)
  );
  sky130_fd_sc_hd__inv_2 _3733_ (
    .A(\g_bit[17].g_word[18].r_bit.Q ),
    .Y(_1397_)
  );
  sky130_fd_sc_hd__or3_2 _3734_ (
    .A(_1397_),
    .B(_0780_),
    .C(_0876_),
    .X(_1398_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3735_ (
    .A1(_1392_),
    .A2(_0868_),
    .B1(_1394_),
    .C1(_1396_),
    .D1(_1398_),
    .Y(_1399_)
  );
  sky130_fd_sc_hd__or4_2 _3736_ (
    .A(_1379_),
    .B(_1381_),
    .C(_1391_),
    .D(_1399_),
    .X(_1400_)
  );
  sky130_fd_sc_hd__or4_2 _3737_ (
    .A(_1365_),
    .B(_1367_),
    .C(_1372_),
    .D(_1400_),
    .X(_1401_)
  );
  sky130_fd_sc_hd__buf_1 _3738_ (
    .A(_1401_),
    .X(\g_bit[17].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _3739_ (
    .A1(\g_bit[17].g_word[30].r_bit.Q ),
    .A2(_0883_),
    .A3(_0884_),
    .B1(_0885_),
    .B2(\g_bit[17].g_word[28].r_bit.Q ),
    .X(_1402_)
  );
  sky130_fd_sc_hd__a221o_2 _3740_ (
    .A1(\g_bit[17].g_word[4].r_bit.Q ),
    .A2(_0881_),
    .B1(_0882_),
    .B2(\g_bit[17].g_word[26].r_bit.Q ),
    .C1(_1402_),
    .X(_1403_)
  );
  sky130_fd_sc_hd__a22o_2 _3741_ (
    .A1(\g_bit[17].g_word[5].r_bit.Q ),
    .A2(_0890_),
    .B1(_0891_),
    .B2(\g_bit[17].g_word[2].r_bit.Q ),
    .X(_1404_)
  );
  sky130_fd_sc_hd__a221o_2 _3742_ (
    .A1(\g_bit[17].g_word[25].r_bit.Q ),
    .A2(_0888_),
    .B1(_0889_),
    .B2(\g_bit[17].g_word[31].r_bit.Q ),
    .C1(_1404_),
    .X(_1405_)
  );
  sky130_fd_sc_hd__a22o_2 _3743_ (
    .A1(\g_bit[17].g_word[13].r_bit.Q ),
    .A2(_0894_),
    .B1(_0895_),
    .B2(\g_bit[17].g_word[15].r_bit.Q ),
    .X(_1406_)
  );
  sky130_fd_sc_hd__a22o_2 _3744_ (
    .A1(\g_bit[17].g_word[20].r_bit.Q ),
    .A2(_0897_),
    .B1(_0898_),
    .B2(\g_bit[17].g_word[11].r_bit.Q ),
    .X(_1407_)
  );
  sky130_fd_sc_hd__a22o_2 _3745_ (
    .A1(\g_bit[17].g_word[19].r_bit.Q ),
    .A2(_0900_),
    .B1(_0901_),
    .B2(\g_bit[17].g_word[21].r_bit.Q ),
    .X(_1408_)
  );
  sky130_fd_sc_hd__a22o_2 _3746_ (
    .A1(\g_bit[17].g_word[17].r_bit.Q ),
    .A2(_0903_),
    .B1(_0904_),
    .B2(\g_bit[17].g_word[12].r_bit.Q ),
    .X(_1409_)
  );
  sky130_fd_sc_hd__or4_2 _3747_ (
    .A(_1406_),
    .B(_1407_),
    .C(_1408_),
    .D(_1409_),
    .X(_1410_)
  );
  sky130_fd_sc_hd__buf_1 _3748_ (
    .A(_0209_),
    .X(_1411_)
  );
  sky130_fd_sc_hd__nor3_2 _3749_ (
    .A(_1373_),
    .B(_0794_),
    .C(_1411_),
    .Y(_1412_)
  );
  sky130_fd_sc_hd__nor3_2 _3750_ (
    .A(_1376_),
    .B(_0909_),
    .C(_0796_),
    .Y(_1413_)
  );
  sky130_fd_sc_hd__and3_2 _3751_ (
    .A(\g_bit[17].g_word[24].r_bit.Q ),
    .B(_0983_),
    .C(_0798_),
    .X(_1414_)
  );
  sky130_fd_sc_hd__a2111o_2 _3752_ (
    .A1(\g_bit[17].g_word[29].r_bit.Q ),
    .A2(_0907_),
    .B1(_1412_),
    .C1(_1413_),
    .D1(_1414_),
    .X(_1415_)
  );
  sky130_fd_sc_hd__and3_2 _3753_ (
    .A(\g_bit[17].g_word[27].r_bit.Q ),
    .B(_0915_),
    .C(_0916_),
    .X(_1416_)
  );
  sky130_fd_sc_hd__a221o_2 _3754_ (
    .A1(\g_bit[17].g_word[6].r_bit.Q ),
    .A2(_0913_),
    .B1(_0914_),
    .B2(\g_bit[17].g_word[1].r_bit.Q ),
    .C1(_1416_),
    .X(_1417_)
  );
  sky130_fd_sc_hd__buf_1 _3755_ (
    .A(_0177_),
    .X(_1418_)
  );
  sky130_fd_sc_hd__or3_2 _3756_ (
    .A(_1383_),
    .B(_1169_),
    .C(_1418_),
    .X(_1419_)
  );
  sky130_fd_sc_hd__or3_2 _3757_ (
    .A(_1386_),
    .B(_1293_),
    .C(_0921_),
    .X(_1420_)
  );
  sky130_fd_sc_hd__buf_1 _3758_ (
    .A(_0144_),
    .X(_1421_)
  );
  sky130_fd_sc_hd__or3_2 _3759_ (
    .A(_1388_),
    .B(_1421_),
    .C(_0923_),
    .X(_1422_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3760_ (
    .A1(_1382_),
    .A2(_0919_),
    .B1(_1419_),
    .C1(_1420_),
    .D1(_1422_),
    .Y(_1423_)
  );
  sky130_fd_sc_hd__or3_2 _3761_ (
    .A(_1393_),
    .B(_0927_),
    .C(_1357_),
    .X(_1424_)
  );
  sky130_fd_sc_hd__or3_2 _3762_ (
    .A(_1395_),
    .B(_0929_),
    .C(_0808_),
    .X(_1425_)
  );
  sky130_fd_sc_hd__or3_2 _3763_ (
    .A(_1397_),
    .B(_0810_),
    .C(_0931_),
    .X(_1426_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3764_ (
    .A1(_1392_),
    .A2(_0926_),
    .B1(_1424_),
    .C1(_1425_),
    .D1(_1426_),
    .Y(_1427_)
  );
  sky130_fd_sc_hd__or4_2 _3765_ (
    .A(_1415_),
    .B(_1417_),
    .C(_1423_),
    .D(_1427_),
    .X(_1428_)
  );
  sky130_fd_sc_hd__or4_2 _3766_ (
    .A(_1403_),
    .B(_1405_),
    .C(_1410_),
    .D(_1428_),
    .X(_1429_)
  );
  sky130_fd_sc_hd__buf_1 _3767_ (
    .A(_1429_),
    .X(\g_bit[17].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _3768_ (
    .A1(\g_bit[18].g_word[30].r_bit.Q ),
    .A2(_0817_),
    .A3(_0818_),
    .B1(_0819_),
    .B2(\g_bit[18].g_word[28].r_bit.Q ),
    .X(_1430_)
  );
  sky130_fd_sc_hd__a221o_2 _3769_ (
    .A1(\g_bit[18].g_word[4].r_bit.Q ),
    .A2(_0815_),
    .B1(_0816_),
    .B2(\g_bit[18].g_word[26].r_bit.Q ),
    .C1(_1430_),
    .X(_1431_)
  );
  sky130_fd_sc_hd__a22o_2 _3770_ (
    .A1(\g_bit[18].g_word[5].r_bit.Q ),
    .A2(_0824_),
    .B1(_0825_),
    .B2(\g_bit[18].g_word[2].r_bit.Q ),
    .X(_1432_)
  );
  sky130_fd_sc_hd__a221o_2 _3771_ (
    .A1(\g_bit[18].g_word[25].r_bit.Q ),
    .A2(_0822_),
    .B1(_0823_),
    .B2(\g_bit[18].g_word[31].r_bit.Q ),
    .C1(_1432_),
    .X(_1433_)
  );
  sky130_fd_sc_hd__a22o_2 _3772_ (
    .A1(\g_bit[18].g_word[13].r_bit.Q ),
    .A2(_0828_),
    .B1(_0829_),
    .B2(\g_bit[18].g_word[15].r_bit.Q ),
    .X(_1434_)
  );
  sky130_fd_sc_hd__a22o_2 _3773_ (
    .A1(\g_bit[18].g_word[11].r_bit.Q ),
    .A2(_0831_),
    .B1(_0832_),
    .B2(\g_bit[18].g_word[20].r_bit.Q ),
    .X(_1435_)
  );
  sky130_fd_sc_hd__a22o_2 _3774_ (
    .A1(\g_bit[18].g_word[19].r_bit.Q ),
    .A2(_0834_),
    .B1(_0835_),
    .B2(\g_bit[18].g_word[21].r_bit.Q ),
    .X(_1436_)
  );
  sky130_fd_sc_hd__a22o_2 _3775_ (
    .A1(\g_bit[18].g_word[17].r_bit.Q ),
    .A2(_0837_),
    .B1(_0838_),
    .B2(\g_bit[18].g_word[12].r_bit.Q ),
    .X(_1437_)
  );
  sky130_fd_sc_hd__or4_2 _3776_ (
    .A(_1434_),
    .B(_1435_),
    .C(_1436_),
    .D(_1437_),
    .X(_1438_)
  );
  sky130_fd_sc_hd__inv_2 _3777_ (
    .A(\g_bit[18].g_word[7].r_bit.Q ),
    .Y(_1439_)
  );
  sky130_fd_sc_hd__buf_1 _3778_ (
    .A(_0003_),
    .X(_1440_)
  );
  sky130_fd_sc_hd__nor3_2 _3779_ (
    .A(_1439_),
    .B(_1374_),
    .C(_1440_),
    .Y(_1441_)
  );
  sky130_fd_sc_hd__inv_2 _3780_ (
    .A(\g_bit[18].g_word[3].r_bit.Q ),
    .Y(_1442_)
  );
  sky130_fd_sc_hd__nor3_2 _3781_ (
    .A(_1442_),
    .B(_0845_),
    .C(_0846_),
    .Y(_1443_)
  );
  sky130_fd_sc_hd__buf_1 _3782_ (
    .A(_0077_),
    .X(_1444_)
  );
  sky130_fd_sc_hd__and3_2 _3783_ (
    .A(\g_bit[18].g_word[24].r_bit.Q ),
    .B(_1444_),
    .C(_0949_),
    .X(_1445_)
  );
  sky130_fd_sc_hd__a2111o_2 _3784_ (
    .A1(\g_bit[18].g_word[29].r_bit.Q ),
    .A2(_0841_),
    .B1(_1441_),
    .C1(_1443_),
    .D1(_1445_),
    .X(_1446_)
  );
  sky130_fd_sc_hd__and3_2 _3785_ (
    .A(\g_bit[18].g_word[27].r_bit.Q ),
    .B(_0852_),
    .C(_0853_),
    .X(_1447_)
  );
  sky130_fd_sc_hd__a221o_2 _3786_ (
    .A1(\g_bit[18].g_word[6].r_bit.Q ),
    .A2(_0850_),
    .B1(_0851_),
    .B2(\g_bit[18].g_word[1].r_bit.Q ),
    .C1(_1447_),
    .X(_1448_)
  );
  sky130_fd_sc_hd__inv_2 _3787_ (
    .A(\g_bit[18].g_word[23].r_bit.Q ),
    .Y(_1449_)
  );
  sky130_fd_sc_hd__inv_2 _3788_ (
    .A(\g_bit[18].g_word[10].r_bit.Q ),
    .Y(_1450_)
  );
  sky130_fd_sc_hd__or3_2 _3789_ (
    .A(_1450_),
    .B(_1137_),
    .C(_1384_),
    .X(_1451_)
  );
  sky130_fd_sc_hd__inv_2 _3790_ (
    .A(\g_bit[18].g_word[9].r_bit.Q ),
    .Y(_1452_)
  );
  sky130_fd_sc_hd__or3_2 _3791_ (
    .A(_1452_),
    .B(_1261_),
    .C(_0861_),
    .X(_1453_)
  );
  sky130_fd_sc_hd__inv_2 _3792_ (
    .A(\g_bit[18].g_word[8].r_bit.Q ),
    .Y(_1454_)
  );
  sky130_fd_sc_hd__or3_2 _3793_ (
    .A(_1454_),
    .B(_1389_),
    .C(_0864_),
    .X(_1455_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3794_ (
    .A1(_1449_),
    .A2(_0857_),
    .B1(_1451_),
    .C1(_1453_),
    .D1(_1455_),
    .Y(_1456_)
  );
  sky130_fd_sc_hd__inv_2 _3795_ (
    .A(\g_bit[18].g_word[22].r_bit.Q ),
    .Y(_1457_)
  );
  sky130_fd_sc_hd__inv_2 _3796_ (
    .A(\g_bit[18].g_word[16].r_bit.Q ),
    .Y(_1458_)
  );
  sky130_fd_sc_hd__or3_2 _3797_ (
    .A(_1458_),
    .B(_1268_),
    .C(_0870_),
    .X(_1459_)
  );
  sky130_fd_sc_hd__inv_2 _3798_ (
    .A(\g_bit[18].g_word[14].r_bit.Q ),
    .Y(_1460_)
  );
  sky130_fd_sc_hd__buf_1 _3799_ (
    .A(_0028_),
    .X(_1461_)
  );
  sky130_fd_sc_hd__or3_2 _3800_ (
    .A(_1460_),
    .B(_0873_),
    .C(_1461_),
    .X(_1462_)
  );
  sky130_fd_sc_hd__inv_2 _3801_ (
    .A(\g_bit[18].g_word[18].r_bit.Q ),
    .Y(_1463_)
  );
  sky130_fd_sc_hd__buf_1 _3802_ (
    .A(_0046_),
    .X(_1464_)
  );
  sky130_fd_sc_hd__or3_2 _3803_ (
    .A(_1463_),
    .B(_1464_),
    .C(_0876_),
    .X(_1465_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3804_ (
    .A1(_1457_),
    .A2(_0868_),
    .B1(_1459_),
    .C1(_1462_),
    .D1(_1465_),
    .Y(_1466_)
  );
  sky130_fd_sc_hd__or4_2 _3805_ (
    .A(_1446_),
    .B(_1448_),
    .C(_1456_),
    .D(_1466_),
    .X(_1467_)
  );
  sky130_fd_sc_hd__or4_2 _3806_ (
    .A(_1431_),
    .B(_1433_),
    .C(_1438_),
    .D(_1467_),
    .X(_1468_)
  );
  sky130_fd_sc_hd__buf_1 _3807_ (
    .A(_1468_),
    .X(\g_bit[18].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _3808_ (
    .A1(\g_bit[18].g_word[30].r_bit.Q ),
    .A2(_0883_),
    .A3(_0884_),
    .B1(_0885_),
    .B2(\g_bit[18].g_word[28].r_bit.Q ),
    .X(_1469_)
  );
  sky130_fd_sc_hd__a221o_2 _3809_ (
    .A1(\g_bit[18].g_word[4].r_bit.Q ),
    .A2(_0881_),
    .B1(_0882_),
    .B2(\g_bit[18].g_word[26].r_bit.Q ),
    .C1(_1469_),
    .X(_1470_)
  );
  sky130_fd_sc_hd__a22o_2 _3810_ (
    .A1(\g_bit[18].g_word[5].r_bit.Q ),
    .A2(_0890_),
    .B1(_0891_),
    .B2(\g_bit[18].g_word[2].r_bit.Q ),
    .X(_1471_)
  );
  sky130_fd_sc_hd__a221o_2 _3811_ (
    .A1(\g_bit[18].g_word[25].r_bit.Q ),
    .A2(_0888_),
    .B1(_0889_),
    .B2(\g_bit[18].g_word[31].r_bit.Q ),
    .C1(_1471_),
    .X(_1472_)
  );
  sky130_fd_sc_hd__a22o_2 _3812_ (
    .A1(\g_bit[18].g_word[13].r_bit.Q ),
    .A2(_0894_),
    .B1(_0895_),
    .B2(\g_bit[18].g_word[15].r_bit.Q ),
    .X(_1473_)
  );
  sky130_fd_sc_hd__a22o_2 _3813_ (
    .A1(\g_bit[18].g_word[20].r_bit.Q ),
    .A2(_0897_),
    .B1(_0898_),
    .B2(\g_bit[18].g_word[11].r_bit.Q ),
    .X(_1474_)
  );
  sky130_fd_sc_hd__a22o_2 _3814_ (
    .A1(\g_bit[18].g_word[19].r_bit.Q ),
    .A2(_0900_),
    .B1(_0901_),
    .B2(\g_bit[18].g_word[21].r_bit.Q ),
    .X(_1475_)
  );
  sky130_fd_sc_hd__a22o_2 _3815_ (
    .A1(\g_bit[18].g_word[17].r_bit.Q ),
    .A2(_0903_),
    .B1(_0904_),
    .B2(\g_bit[18].g_word[12].r_bit.Q ),
    .X(_1476_)
  );
  sky130_fd_sc_hd__or4_2 _3816_ (
    .A(_1473_),
    .B(_1474_),
    .C(_1475_),
    .D(_1476_),
    .X(_1477_)
  );
  sky130_fd_sc_hd__buf_1 _3817_ (
    .A(_0132_),
    .X(_1478_)
  );
  sky130_fd_sc_hd__nor3_2 _3818_ (
    .A(_1439_),
    .B(_1478_),
    .C(_1411_),
    .Y(_1479_)
  );
  sky130_fd_sc_hd__buf_1 _3819_ (
    .A(_0209_),
    .X(_1480_)
  );
  sky130_fd_sc_hd__nor3_2 _3820_ (
    .A(_1442_),
    .B(_0909_),
    .C(_1480_),
    .Y(_1481_)
  );
  sky130_fd_sc_hd__buf_1 _3821_ (
    .A(_0207_),
    .X(_1482_)
  );
  sky130_fd_sc_hd__and3_2 _3822_ (
    .A(\g_bit[18].g_word[24].r_bit.Q ),
    .B(_0983_),
    .C(_1482_),
    .X(_1483_)
  );
  sky130_fd_sc_hd__a2111o_2 _3823_ (
    .A1(\g_bit[18].g_word[29].r_bit.Q ),
    .A2(_0907_),
    .B1(_1479_),
    .C1(_1481_),
    .D1(_1483_),
    .X(_1484_)
  );
  sky130_fd_sc_hd__and3_2 _3824_ (
    .A(\g_bit[18].g_word[27].r_bit.Q ),
    .B(_0915_),
    .C(_0916_),
    .X(_1485_)
  );
  sky130_fd_sc_hd__a221o_2 _3825_ (
    .A1(\g_bit[18].g_word[6].r_bit.Q ),
    .A2(_0913_),
    .B1(_0914_),
    .B2(\g_bit[18].g_word[1].r_bit.Q ),
    .C1(_1485_),
    .X(_1486_)
  );
  sky130_fd_sc_hd__or3_2 _3826_ (
    .A(_1450_),
    .B(_1169_),
    .C(_1418_),
    .X(_1487_)
  );
  sky130_fd_sc_hd__or3_2 _3827_ (
    .A(_1452_),
    .B(_1293_),
    .C(_0921_),
    .X(_1488_)
  );
  sky130_fd_sc_hd__or3_2 _3828_ (
    .A(_1454_),
    .B(_1421_),
    .C(_0923_),
    .X(_1489_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3829_ (
    .A1(_1449_),
    .A2(_0919_),
    .B1(_1487_),
    .C1(_1488_),
    .D1(_1489_),
    .Y(_1490_)
  );
  sky130_fd_sc_hd__or3_2 _3830_ (
    .A(_1458_),
    .B(_0927_),
    .C(_1357_),
    .X(_1491_)
  );
  sky130_fd_sc_hd__buf_1 _3831_ (
    .A(_0157_),
    .X(_1492_)
  );
  sky130_fd_sc_hd__or3_2 _3832_ (
    .A(_1460_),
    .B(_0929_),
    .C(_1492_),
    .X(_1493_)
  );
  sky130_fd_sc_hd__buf_1 _3833_ (
    .A(_0175_),
    .X(_1494_)
  );
  sky130_fd_sc_hd__or3_2 _3834_ (
    .A(_1463_),
    .B(_1494_),
    .C(_0931_),
    .X(_1495_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3835_ (
    .A1(_1457_),
    .A2(_0926_),
    .B1(_1491_),
    .C1(_1493_),
    .D1(_1495_),
    .Y(_1496_)
  );
  sky130_fd_sc_hd__or4_2 _3836_ (
    .A(_1484_),
    .B(_1486_),
    .C(_1490_),
    .D(_1496_),
    .X(_1497_)
  );
  sky130_fd_sc_hd__or4_2 _3837_ (
    .A(_1470_),
    .B(_1472_),
    .C(_1477_),
    .D(_1497_),
    .X(_1498_)
  );
  sky130_fd_sc_hd__buf_1 _3838_ (
    .A(_1498_),
    .X(\g_bit[18].r_rs2.D )
  );
  sky130_fd_sc_hd__buf_1 _3839_ (
    .A(_0013_),
    .X(_1499_)
  );
  sky130_fd_sc_hd__buf_1 _3840_ (
    .A(_0020_),
    .X(_1500_)
  );
  sky130_fd_sc_hd__buf_1 _3841_ (
    .A(_0022_),
    .X(_1501_)
  );
  sky130_fd_sc_hd__buf_1 _3842_ (
    .A(_0024_),
    .X(_1502_)
  );
  sky130_fd_sc_hd__buf_1 _3843_ (
    .A(_0029_),
    .X(_1503_)
  );
  sky130_fd_sc_hd__a32o_2 _3844_ (
    .A1(\g_bit[19].g_word[30].r_bit.Q ),
    .A2(_1501_),
    .A3(_1502_),
    .B1(_1503_),
    .B2(\g_bit[19].g_word[28].r_bit.Q ),
    .X(_1504_)
  );
  sky130_fd_sc_hd__a221o_2 _3845_ (
    .A1(\g_bit[19].g_word[4].r_bit.Q ),
    .A2(_1499_),
    .B1(_1500_),
    .B2(\g_bit[19].g_word[26].r_bit.Q ),
    .C1(_1504_),
    .X(_1505_)
  );
  sky130_fd_sc_hd__buf_1 _3846_ (
    .A(_0034_),
    .X(_1506_)
  );
  sky130_fd_sc_hd__buf_1 _3847_ (
    .A(_0038_),
    .X(_1507_)
  );
  sky130_fd_sc_hd__buf_1 _3848_ (
    .A(_0042_),
    .X(_1508_)
  );
  sky130_fd_sc_hd__buf_1 _3849_ (
    .A(_0049_),
    .X(_1509_)
  );
  sky130_fd_sc_hd__a22o_2 _3850_ (
    .A1(\g_bit[19].g_word[5].r_bit.Q ),
    .A2(_1508_),
    .B1(_1509_),
    .B2(\g_bit[19].g_word[2].r_bit.Q ),
    .X(_1510_)
  );
  sky130_fd_sc_hd__a221o_2 _3851_ (
    .A1(\g_bit[19].g_word[25].r_bit.Q ),
    .A2(_1506_),
    .B1(_1507_),
    .B2(\g_bit[19].g_word[31].r_bit.Q ),
    .C1(_1510_),
    .X(_1511_)
  );
  sky130_fd_sc_hd__buf_1 _3852_ (
    .A(_0053_),
    .X(_1512_)
  );
  sky130_fd_sc_hd__buf_1 _3853_ (
    .A(_0056_),
    .X(_1513_)
  );
  sky130_fd_sc_hd__a22o_2 _3854_ (
    .A1(\g_bit[19].g_word[13].r_bit.Q ),
    .A2(_1512_),
    .B1(_1513_),
    .B2(\g_bit[19].g_word[15].r_bit.Q ),
    .X(_1514_)
  );
  sky130_fd_sc_hd__buf_1 _3855_ (
    .A(_0059_),
    .X(_1515_)
  );
  sky130_fd_sc_hd__buf_1 _3856_ (
    .A(_0061_),
    .X(_1516_)
  );
  sky130_fd_sc_hd__a22o_2 _3857_ (
    .A1(\g_bit[19].g_word[11].r_bit.Q ),
    .A2(_1515_),
    .B1(_1516_),
    .B2(\g_bit[19].g_word[20].r_bit.Q ),
    .X(_1517_)
  );
  sky130_fd_sc_hd__buf_1 _3858_ (
    .A(_0064_),
    .X(_1518_)
  );
  sky130_fd_sc_hd__buf_1 _3859_ (
    .A(_0066_),
    .X(_1519_)
  );
  sky130_fd_sc_hd__a22o_2 _3860_ (
    .A1(\g_bit[19].g_word[19].r_bit.Q ),
    .A2(_1518_),
    .B1(_1519_),
    .B2(\g_bit[19].g_word[21].r_bit.Q ),
    .X(_1520_)
  );
  sky130_fd_sc_hd__buf_1 _3861_ (
    .A(_0069_),
    .X(_1521_)
  );
  sky130_fd_sc_hd__buf_1 _3862_ (
    .A(_0071_),
    .X(_1522_)
  );
  sky130_fd_sc_hd__a22o_2 _3863_ (
    .A1(\g_bit[19].g_word[17].r_bit.Q ),
    .A2(_1521_),
    .B1(_1522_),
    .B2(\g_bit[19].g_word[12].r_bit.Q ),
    .X(_1523_)
  );
  sky130_fd_sc_hd__or4_2 _3864_ (
    .A(_1514_),
    .B(_1517_),
    .C(_1520_),
    .D(_1523_),
    .X(_1524_)
  );
  sky130_fd_sc_hd__buf_1 _3865_ (
    .A(_0075_),
    .X(_1525_)
  );
  sky130_fd_sc_hd__inv_2 _3866_ (
    .A(\g_bit[19].g_word[7].r_bit.Q ),
    .Y(_1526_)
  );
  sky130_fd_sc_hd__nor3_2 _3867_ (
    .A(_1526_),
    .B(_1374_),
    .C(_1440_),
    .Y(_1527_)
  );
  sky130_fd_sc_hd__inv_2 _3868_ (
    .A(\g_bit[19].g_word[3].r_bit.Q ),
    .Y(_1528_)
  );
  sky130_fd_sc_hd__buf_1 _3869_ (
    .A(_0045_),
    .X(_1529_)
  );
  sky130_fd_sc_hd__buf_1 _3870_ (
    .A(_0081_),
    .X(_1530_)
  );
  sky130_fd_sc_hd__nor3_2 _3871_ (
    .A(_1528_),
    .B(_1529_),
    .C(_1530_),
    .Y(_1531_)
  );
  sky130_fd_sc_hd__and3_2 _3872_ (
    .A(\g_bit[19].g_word[24].r_bit.Q ),
    .B(_1444_),
    .C(_0949_),
    .X(_1532_)
  );
  sky130_fd_sc_hd__a2111o_2 _3873_ (
    .A1(\g_bit[19].g_word[29].r_bit.Q ),
    .A2(_1525_),
    .B1(_1527_),
    .C1(_1531_),
    .D1(_1532_),
    .X(_1533_)
  );
  sky130_fd_sc_hd__buf_1 _3874_ (
    .A(_0089_),
    .X(_1534_)
  );
  sky130_fd_sc_hd__buf_1 _3875_ (
    .A(_0091_),
    .X(_1535_)
  );
  sky130_fd_sc_hd__buf_1 _3876_ (
    .A(_0093_),
    .X(_1536_)
  );
  sky130_fd_sc_hd__buf_1 _3877_ (
    .A(_0077_),
    .X(_1537_)
  );
  sky130_fd_sc_hd__and3_2 _3878_ (
    .A(\g_bit[19].g_word[27].r_bit.Q ),
    .B(_1536_),
    .C(_1537_),
    .X(_1538_)
  );
  sky130_fd_sc_hd__a221o_2 _3879_ (
    .A1(\g_bit[19].g_word[6].r_bit.Q ),
    .A2(_1534_),
    .B1(_1535_),
    .B2(\g_bit[19].g_word[1].r_bit.Q ),
    .C1(_1538_),
    .X(_1539_)
  );
  sky130_fd_sc_hd__inv_2 _3880_ (
    .A(\g_bit[19].g_word[23].r_bit.Q ),
    .Y(_1540_)
  );
  sky130_fd_sc_hd__buf_1 _3881_ (
    .A(_0100_),
    .X(_1541_)
  );
  sky130_fd_sc_hd__inv_2 _3882_ (
    .A(\g_bit[19].g_word[10].r_bit.Q ),
    .Y(_1542_)
  );
  sky130_fd_sc_hd__or3_2 _3883_ (
    .A(_1542_),
    .B(_1137_),
    .C(_1384_),
    .X(_1543_)
  );
  sky130_fd_sc_hd__inv_2 _3884_ (
    .A(\g_bit[19].g_word[9].r_bit.Q ),
    .Y(_1544_)
  );
  sky130_fd_sc_hd__buf_1 _3885_ (
    .A(_0041_),
    .X(_1545_)
  );
  sky130_fd_sc_hd__or3_2 _3886_ (
    .A(_1544_),
    .B(_1261_),
    .C(_1545_),
    .X(_1546_)
  );
  sky130_fd_sc_hd__inv_2 _3887_ (
    .A(\g_bit[19].g_word[8].r_bit.Q ),
    .Y(_1547_)
  );
  sky130_fd_sc_hd__buf_1 _3888_ (
    .A(_0011_),
    .X(_1548_)
  );
  sky130_fd_sc_hd__or3_2 _3889_ (
    .A(_1547_),
    .B(_1389_),
    .C(_1548_),
    .X(_1549_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3890_ (
    .A1(_1540_),
    .A2(_1541_),
    .B1(_1543_),
    .C1(_1546_),
    .D1(_1549_),
    .Y(_1550_)
  );
  sky130_fd_sc_hd__inv_2 _3891_ (
    .A(\g_bit[19].g_word[22].r_bit.Q ),
    .Y(_1551_)
  );
  sky130_fd_sc_hd__buf_1 _3892_ (
    .A(_0115_),
    .X(_1552_)
  );
  sky130_fd_sc_hd__inv_2 _3893_ (
    .A(\g_bit[19].g_word[16].r_bit.Q ),
    .Y(_1553_)
  );
  sky130_fd_sc_hd__buf_1 _3894_ (
    .A(_0026_),
    .X(_1554_)
  );
  sky130_fd_sc_hd__or3_2 _3895_ (
    .A(_1553_),
    .B(_1268_),
    .C(_1554_),
    .X(_1555_)
  );
  sky130_fd_sc_hd__inv_2 _3896_ (
    .A(\g_bit[19].g_word[14].r_bit.Q ),
    .Y(_1556_)
  );
  sky130_fd_sc_hd__buf_1 _3897_ (
    .A(_0048_),
    .X(_1557_)
  );
  sky130_fd_sc_hd__or3_2 _3898_ (
    .A(_1556_),
    .B(_1557_),
    .C(_1461_),
    .X(_1558_)
  );
  sky130_fd_sc_hd__inv_2 _3899_ (
    .A(\g_bit[19].g_word[18].r_bit.Q ),
    .Y(_1559_)
  );
  sky130_fd_sc_hd__buf_1 _3900_ (
    .A(_0018_),
    .X(_1560_)
  );
  sky130_fd_sc_hd__or3_2 _3901_ (
    .A(_1559_),
    .B(_1464_),
    .C(_1560_),
    .X(_1561_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3902_ (
    .A1(_1551_),
    .A2(_1552_),
    .B1(_1555_),
    .C1(_1558_),
    .D1(_1561_),
    .Y(_1562_)
  );
  sky130_fd_sc_hd__or4_2 _3903_ (
    .A(_1533_),
    .B(_1539_),
    .C(_1550_),
    .D(_1562_),
    .X(_1563_)
  );
  sky130_fd_sc_hd__or4_2 _3904_ (
    .A(_1505_),
    .B(_1511_),
    .C(_1524_),
    .D(_1563_),
    .X(_1564_)
  );
  sky130_fd_sc_hd__buf_1 _3905_ (
    .A(_1564_),
    .X(\g_bit[19].r_rs1.D )
  );
  sky130_fd_sc_hd__buf_1 _3906_ (
    .A(_0142_),
    .X(_1565_)
  );
  sky130_fd_sc_hd__buf_1 _3907_ (
    .A(_0149_),
    .X(_1566_)
  );
  sky130_fd_sc_hd__buf_1 _3908_ (
    .A(_0151_),
    .X(_1567_)
  );
  sky130_fd_sc_hd__buf_1 _3909_ (
    .A(_0153_),
    .X(_1568_)
  );
  sky130_fd_sc_hd__buf_1 _3910_ (
    .A(_0158_),
    .X(_1569_)
  );
  sky130_fd_sc_hd__a32o_2 _3911_ (
    .A1(\g_bit[19].g_word[30].r_bit.Q ),
    .A2(_1567_),
    .A3(_1568_),
    .B1(_1569_),
    .B2(\g_bit[19].g_word[28].r_bit.Q ),
    .X(_1570_)
  );
  sky130_fd_sc_hd__a221o_2 _3912_ (
    .A1(\g_bit[19].g_word[4].r_bit.Q ),
    .A2(_1565_),
    .B1(_1566_),
    .B2(\g_bit[19].g_word[26].r_bit.Q ),
    .C1(_1570_),
    .X(_1571_)
  );
  sky130_fd_sc_hd__buf_1 _3913_ (
    .A(_0163_),
    .X(_1572_)
  );
  sky130_fd_sc_hd__buf_1 _3914_ (
    .A(_0167_),
    .X(_1573_)
  );
  sky130_fd_sc_hd__buf_1 _3915_ (
    .A(_0171_),
    .X(_1574_)
  );
  sky130_fd_sc_hd__buf_1 _3916_ (
    .A(_0178_),
    .X(_1575_)
  );
  sky130_fd_sc_hd__a22o_2 _3917_ (
    .A1(\g_bit[19].g_word[5].r_bit.Q ),
    .A2(_1574_),
    .B1(_1575_),
    .B2(\g_bit[19].g_word[2].r_bit.Q ),
    .X(_1576_)
  );
  sky130_fd_sc_hd__a221o_2 _3918_ (
    .A1(\g_bit[19].g_word[25].r_bit.Q ),
    .A2(_1572_),
    .B1(_1573_),
    .B2(\g_bit[19].g_word[31].r_bit.Q ),
    .C1(_1576_),
    .X(_1577_)
  );
  sky130_fd_sc_hd__buf_1 _3919_ (
    .A(_0182_),
    .X(_1578_)
  );
  sky130_fd_sc_hd__buf_1 _3920_ (
    .A(_0185_),
    .X(_1579_)
  );
  sky130_fd_sc_hd__a22o_2 _3921_ (
    .A1(\g_bit[19].g_word[13].r_bit.Q ),
    .A2(_1578_),
    .B1(_1579_),
    .B2(\g_bit[19].g_word[15].r_bit.Q ),
    .X(_1580_)
  );
  sky130_fd_sc_hd__buf_1 _3922_ (
    .A(_0188_),
    .X(_1581_)
  );
  sky130_fd_sc_hd__buf_1 _3923_ (
    .A(_0190_),
    .X(_1582_)
  );
  sky130_fd_sc_hd__a22o_2 _3924_ (
    .A1(\g_bit[19].g_word[20].r_bit.Q ),
    .A2(_1581_),
    .B1(_1582_),
    .B2(\g_bit[19].g_word[11].r_bit.Q ),
    .X(_1583_)
  );
  sky130_fd_sc_hd__buf_1 _3925_ (
    .A(_0193_),
    .X(_1584_)
  );
  sky130_fd_sc_hd__buf_1 _3926_ (
    .A(_0195_),
    .X(_1585_)
  );
  sky130_fd_sc_hd__a22o_2 _3927_ (
    .A1(\g_bit[19].g_word[19].r_bit.Q ),
    .A2(_1584_),
    .B1(_1585_),
    .B2(\g_bit[19].g_word[21].r_bit.Q ),
    .X(_1586_)
  );
  sky130_fd_sc_hd__buf_1 _3928_ (
    .A(_0198_),
    .X(_1587_)
  );
  sky130_fd_sc_hd__buf_1 _3929_ (
    .A(_0200_),
    .X(_1588_)
  );
  sky130_fd_sc_hd__a22o_2 _3930_ (
    .A1(\g_bit[19].g_word[17].r_bit.Q ),
    .A2(_1587_),
    .B1(_1588_),
    .B2(\g_bit[19].g_word[12].r_bit.Q ),
    .X(_1589_)
  );
  sky130_fd_sc_hd__or4_2 _3931_ (
    .A(_1580_),
    .B(_1583_),
    .C(_1586_),
    .D(_1589_),
    .X(_1590_)
  );
  sky130_fd_sc_hd__buf_1 _3932_ (
    .A(_0204_),
    .X(_1591_)
  );
  sky130_fd_sc_hd__nor3_2 _3933_ (
    .A(_1526_),
    .B(_1478_),
    .C(_1411_),
    .Y(_1592_)
  );
  sky130_fd_sc_hd__buf_1 _3934_ (
    .A(_0174_),
    .X(_1593_)
  );
  sky130_fd_sc_hd__nor3_2 _3935_ (
    .A(_1528_),
    .B(_1593_),
    .C(_1480_),
    .Y(_1594_)
  );
  sky130_fd_sc_hd__and3_2 _3936_ (
    .A(\g_bit[19].g_word[24].r_bit.Q ),
    .B(_0983_),
    .C(_1482_),
    .X(_1595_)
  );
  sky130_fd_sc_hd__a2111o_2 _3937_ (
    .A1(\g_bit[19].g_word[29].r_bit.Q ),
    .A2(_1591_),
    .B1(_1592_),
    .C1(_1594_),
    .D1(_1595_),
    .X(_1596_)
  );
  sky130_fd_sc_hd__buf_1 _3938_ (
    .A(_0215_),
    .X(_1597_)
  );
  sky130_fd_sc_hd__buf_1 _3939_ (
    .A(_0217_),
    .X(_1598_)
  );
  sky130_fd_sc_hd__buf_1 _3940_ (
    .A(_0219_),
    .X(_1599_)
  );
  sky130_fd_sc_hd__buf_1 _3941_ (
    .A(_0207_),
    .X(_1600_)
  );
  sky130_fd_sc_hd__and3_2 _3942_ (
    .A(\g_bit[19].g_word[27].r_bit.Q ),
    .B(_1599_),
    .C(_1600_),
    .X(_1601_)
  );
  sky130_fd_sc_hd__a221o_2 _3943_ (
    .A1(\g_bit[19].g_word[6].r_bit.Q ),
    .A2(_1597_),
    .B1(_1598_),
    .B2(\g_bit[19].g_word[1].r_bit.Q ),
    .C1(_1601_),
    .X(_1602_)
  );
  sky130_fd_sc_hd__buf_1 _3944_ (
    .A(_0225_),
    .X(_1603_)
  );
  sky130_fd_sc_hd__or3_2 _3945_ (
    .A(_1542_),
    .B(_1169_),
    .C(_1418_),
    .X(_1604_)
  );
  sky130_fd_sc_hd__buf_1 _3946_ (
    .A(_0170_),
    .X(_1605_)
  );
  sky130_fd_sc_hd__or3_2 _3947_ (
    .A(_1544_),
    .B(_1293_),
    .C(_1605_),
    .X(_1606_)
  );
  sky130_fd_sc_hd__buf_1 _3948_ (
    .A(_0140_),
    .X(_1607_)
  );
  sky130_fd_sc_hd__or3_2 _3949_ (
    .A(_1547_),
    .B(_1421_),
    .C(_1607_),
    .X(_1608_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3950_ (
    .A1(_1540_),
    .A2(_1603_),
    .B1(_1604_),
    .C1(_1606_),
    .D1(_1608_),
    .Y(_1609_)
  );
  sky130_fd_sc_hd__buf_1 _3951_ (
    .A(_0236_),
    .X(_1610_)
  );
  sky130_fd_sc_hd__buf_1 _3952_ (
    .A(_0155_),
    .X(_1611_)
  );
  sky130_fd_sc_hd__or3_2 _3953_ (
    .A(_1553_),
    .B(_1611_),
    .C(_1357_),
    .X(_1612_)
  );
  sky130_fd_sc_hd__buf_1 _3954_ (
    .A(_0177_),
    .X(_1613_)
  );
  sky130_fd_sc_hd__or3_2 _3955_ (
    .A(_1556_),
    .B(_1613_),
    .C(_1492_),
    .X(_1614_)
  );
  sky130_fd_sc_hd__buf_1 _3956_ (
    .A(_0147_),
    .X(_1615_)
  );
  sky130_fd_sc_hd__or3_2 _3957_ (
    .A(_1559_),
    .B(_1494_),
    .C(_1615_),
    .X(_1616_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3958_ (
    .A1(_1551_),
    .A2(_1610_),
    .B1(_1612_),
    .C1(_1614_),
    .D1(_1616_),
    .Y(_1617_)
  );
  sky130_fd_sc_hd__or4_2 _3959_ (
    .A(_1596_),
    .B(_1602_),
    .C(_1609_),
    .D(_1617_),
    .X(_1618_)
  );
  sky130_fd_sc_hd__or4_2 _3960_ (
    .A(_1571_),
    .B(_1577_),
    .C(_1590_),
    .D(_1618_),
    .X(_1619_)
  );
  sky130_fd_sc_hd__buf_1 _3961_ (
    .A(_1619_),
    .X(\g_bit[19].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _3962_ (
    .A1(\g_bit[20].g_word[30].r_bit.Q ),
    .A2(_1501_),
    .A3(_1502_),
    .B1(_1503_),
    .B2(\g_bit[20].g_word[28].r_bit.Q ),
    .X(_1620_)
  );
  sky130_fd_sc_hd__a221o_2 _3963_ (
    .A1(\g_bit[20].g_word[4].r_bit.Q ),
    .A2(_1499_),
    .B1(_1500_),
    .B2(\g_bit[20].g_word[26].r_bit.Q ),
    .C1(_1620_),
    .X(_1621_)
  );
  sky130_fd_sc_hd__a22o_2 _3964_ (
    .A1(\g_bit[20].g_word[5].r_bit.Q ),
    .A2(_1508_),
    .B1(_1509_),
    .B2(\g_bit[20].g_word[2].r_bit.Q ),
    .X(_1622_)
  );
  sky130_fd_sc_hd__a221o_2 _3965_ (
    .A1(\g_bit[20].g_word[25].r_bit.Q ),
    .A2(_1506_),
    .B1(_1507_),
    .B2(\g_bit[20].g_word[31].r_bit.Q ),
    .C1(_1622_),
    .X(_1623_)
  );
  sky130_fd_sc_hd__a22o_2 _3966_ (
    .A1(\g_bit[20].g_word[13].r_bit.Q ),
    .A2(_1512_),
    .B1(_1513_),
    .B2(\g_bit[20].g_word[15].r_bit.Q ),
    .X(_1624_)
  );
  sky130_fd_sc_hd__a22o_2 _3967_ (
    .A1(\g_bit[20].g_word[11].r_bit.Q ),
    .A2(_1515_),
    .B1(_1516_),
    .B2(\g_bit[20].g_word[20].r_bit.Q ),
    .X(_1625_)
  );
  sky130_fd_sc_hd__a22o_2 _3968_ (
    .A1(\g_bit[20].g_word[19].r_bit.Q ),
    .A2(_1518_),
    .B1(_1519_),
    .B2(\g_bit[20].g_word[21].r_bit.Q ),
    .X(_1626_)
  );
  sky130_fd_sc_hd__a22o_2 _3969_ (
    .A1(\g_bit[20].g_word[17].r_bit.Q ),
    .A2(_1521_),
    .B1(_1522_),
    .B2(\g_bit[20].g_word[12].r_bit.Q ),
    .X(_1627_)
  );
  sky130_fd_sc_hd__or4_2 _3970_ (
    .A(_1624_),
    .B(_1625_),
    .C(_1626_),
    .D(_1627_),
    .X(_1628_)
  );
  sky130_fd_sc_hd__inv_2 _3971_ (
    .A(\g_bit[20].g_word[7].r_bit.Q ),
    .Y(_1629_)
  );
  sky130_fd_sc_hd__nor3_2 _3972_ (
    .A(_1629_),
    .B(_1374_),
    .C(_1440_),
    .Y(_1630_)
  );
  sky130_fd_sc_hd__inv_2 _3973_ (
    .A(\g_bit[20].g_word[3].r_bit.Q ),
    .Y(_1631_)
  );
  sky130_fd_sc_hd__nor3_2 _3974_ (
    .A(_1631_),
    .B(_1529_),
    .C(_1530_),
    .Y(_1632_)
  );
  sky130_fd_sc_hd__buf_1 _3975_ (
    .A(_0078_),
    .X(_1633_)
  );
  sky130_fd_sc_hd__and3_2 _3976_ (
    .A(\g_bit[20].g_word[24].r_bit.Q ),
    .B(_1444_),
    .C(_1633_),
    .X(_1634_)
  );
  sky130_fd_sc_hd__a2111o_2 _3977_ (
    .A1(\g_bit[20].g_word[29].r_bit.Q ),
    .A2(_1525_),
    .B1(_1630_),
    .C1(_1632_),
    .D1(_1634_),
    .X(_1635_)
  );
  sky130_fd_sc_hd__and3_2 _3978_ (
    .A(\g_bit[20].g_word[27].r_bit.Q ),
    .B(_1536_),
    .C(_1537_),
    .X(_1636_)
  );
  sky130_fd_sc_hd__a221o_2 _3979_ (
    .A1(\g_bit[20].g_word[6].r_bit.Q ),
    .A2(_1534_),
    .B1(_1535_),
    .B2(\g_bit[20].g_word[1].r_bit.Q ),
    .C1(_1636_),
    .X(_1637_)
  );
  sky130_fd_sc_hd__inv_2 _3980_ (
    .A(\g_bit[20].g_word[23].r_bit.Q ),
    .Y(_1638_)
  );
  sky130_fd_sc_hd__inv_2 _3981_ (
    .A(\g_bit[20].g_word[10].r_bit.Q ),
    .Y(_1639_)
  );
  sky130_fd_sc_hd__or3_2 _3982_ (
    .A(_1639_),
    .B(_1137_),
    .C(_1384_),
    .X(_1640_)
  );
  sky130_fd_sc_hd__inv_2 _3983_ (
    .A(\g_bit[20].g_word[9].r_bit.Q ),
    .Y(_1641_)
  );
  sky130_fd_sc_hd__or3_2 _3984_ (
    .A(_1641_),
    .B(_1261_),
    .C(_1545_),
    .X(_1642_)
  );
  sky130_fd_sc_hd__inv_2 _3985_ (
    .A(\g_bit[20].g_word[8].r_bit.Q ),
    .Y(_1643_)
  );
  sky130_fd_sc_hd__or3_2 _3986_ (
    .A(_1643_),
    .B(_1389_),
    .C(_1548_),
    .X(_1644_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3987_ (
    .A1(_1638_),
    .A2(_1541_),
    .B1(_1640_),
    .C1(_1642_),
    .D1(_1644_),
    .Y(_1645_)
  );
  sky130_fd_sc_hd__inv_2 _3988_ (
    .A(\g_bit[20].g_word[22].r_bit.Q ),
    .Y(_1646_)
  );
  sky130_fd_sc_hd__inv_2 _3989_ (
    .A(\g_bit[20].g_word[16].r_bit.Q ),
    .Y(_1647_)
  );
  sky130_fd_sc_hd__or3_2 _3990_ (
    .A(_1647_),
    .B(_1268_),
    .C(_1554_),
    .X(_1648_)
  );
  sky130_fd_sc_hd__inv_2 _3991_ (
    .A(\g_bit[20].g_word[14].r_bit.Q ),
    .Y(_1649_)
  );
  sky130_fd_sc_hd__or3_2 _3992_ (
    .A(_1649_),
    .B(_1557_),
    .C(_1461_),
    .X(_1650_)
  );
  sky130_fd_sc_hd__inv_2 _3993_ (
    .A(\g_bit[20].g_word[18].r_bit.Q ),
    .Y(_1651_)
  );
  sky130_fd_sc_hd__or3_2 _3994_ (
    .A(_1651_),
    .B(_1464_),
    .C(_1560_),
    .X(_1652_)
  );
  sky130_fd_sc_hd__o2111ai_2 _3995_ (
    .A1(_1646_),
    .A2(_1552_),
    .B1(_1648_),
    .C1(_1650_),
    .D1(_1652_),
    .Y(_1653_)
  );
  sky130_fd_sc_hd__or4_2 _3996_ (
    .A(_1635_),
    .B(_1637_),
    .C(_1645_),
    .D(_1653_),
    .X(_1654_)
  );
  sky130_fd_sc_hd__or4_2 _3997_ (
    .A(_1621_),
    .B(_1623_),
    .C(_1628_),
    .D(_1654_),
    .X(_1655_)
  );
  sky130_fd_sc_hd__buf_1 _3998_ (
    .A(_1655_),
    .X(\g_bit[20].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _3999_ (
    .A1(\g_bit[20].g_word[30].r_bit.Q ),
    .A2(_1567_),
    .A3(_1568_),
    .B1(_1569_),
    .B2(\g_bit[20].g_word[28].r_bit.Q ),
    .X(_1656_)
  );
  sky130_fd_sc_hd__a221o_2 _4000_ (
    .A1(\g_bit[20].g_word[4].r_bit.Q ),
    .A2(_1565_),
    .B1(_1566_),
    .B2(\g_bit[20].g_word[26].r_bit.Q ),
    .C1(_1656_),
    .X(_1657_)
  );
  sky130_fd_sc_hd__a22o_2 _4001_ (
    .A1(\g_bit[20].g_word[5].r_bit.Q ),
    .A2(_1574_),
    .B1(_1575_),
    .B2(\g_bit[20].g_word[2].r_bit.Q ),
    .X(_1658_)
  );
  sky130_fd_sc_hd__a221o_2 _4002_ (
    .A1(\g_bit[20].g_word[25].r_bit.Q ),
    .A2(_1572_),
    .B1(_1573_),
    .B2(\g_bit[20].g_word[31].r_bit.Q ),
    .C1(_1658_),
    .X(_1659_)
  );
  sky130_fd_sc_hd__a22o_2 _4003_ (
    .A1(\g_bit[20].g_word[13].r_bit.Q ),
    .A2(_1578_),
    .B1(_1579_),
    .B2(\g_bit[20].g_word[15].r_bit.Q ),
    .X(_1660_)
  );
  sky130_fd_sc_hd__a22o_2 _4004_ (
    .A1(\g_bit[20].g_word[20].r_bit.Q ),
    .A2(_1581_),
    .B1(_1582_),
    .B2(\g_bit[20].g_word[11].r_bit.Q ),
    .X(_1661_)
  );
  sky130_fd_sc_hd__a22o_2 _4005_ (
    .A1(\g_bit[20].g_word[19].r_bit.Q ),
    .A2(_1584_),
    .B1(_1585_),
    .B2(\g_bit[20].g_word[21].r_bit.Q ),
    .X(_1662_)
  );
  sky130_fd_sc_hd__a22o_2 _4006_ (
    .A1(\g_bit[20].g_word[17].r_bit.Q ),
    .A2(_1587_),
    .B1(_1588_),
    .B2(\g_bit[20].g_word[12].r_bit.Q ),
    .X(_1663_)
  );
  sky130_fd_sc_hd__or4_2 _4007_ (
    .A(_1660_),
    .B(_1661_),
    .C(_1662_),
    .D(_1663_),
    .X(_1664_)
  );
  sky130_fd_sc_hd__nor3_2 _4008_ (
    .A(_1629_),
    .B(_1478_),
    .C(_1411_),
    .Y(_1665_)
  );
  sky130_fd_sc_hd__nor3_2 _4009_ (
    .A(_1631_),
    .B(_1593_),
    .C(_1480_),
    .Y(_1666_)
  );
  sky130_fd_sc_hd__buf_1 _4010_ (
    .A(_0206_),
    .X(_1667_)
  );
  sky130_fd_sc_hd__and3_2 _4011_ (
    .A(\g_bit[20].g_word[24].r_bit.Q ),
    .B(_1667_),
    .C(_1482_),
    .X(_1668_)
  );
  sky130_fd_sc_hd__a2111o_2 _4012_ (
    .A1(\g_bit[20].g_word[29].r_bit.Q ),
    .A2(_1591_),
    .B1(_1665_),
    .C1(_1666_),
    .D1(_1668_),
    .X(_1669_)
  );
  sky130_fd_sc_hd__and3_2 _4013_ (
    .A(\g_bit[20].g_word[27].r_bit.Q ),
    .B(_1599_),
    .C(_1600_),
    .X(_1670_)
  );
  sky130_fd_sc_hd__a221o_2 _4014_ (
    .A1(\g_bit[20].g_word[6].r_bit.Q ),
    .A2(_1597_),
    .B1(_1598_),
    .B2(\g_bit[20].g_word[1].r_bit.Q ),
    .C1(_1670_),
    .X(_1671_)
  );
  sky130_fd_sc_hd__or3_2 _4015_ (
    .A(_1639_),
    .B(_1169_),
    .C(_1418_),
    .X(_1672_)
  );
  sky130_fd_sc_hd__or3_2 _4016_ (
    .A(_1641_),
    .B(_1293_),
    .C(_1605_),
    .X(_1673_)
  );
  sky130_fd_sc_hd__or3_2 _4017_ (
    .A(_1643_),
    .B(_1421_),
    .C(_1607_),
    .X(_1674_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4018_ (
    .A1(_1638_),
    .A2(_1603_),
    .B1(_1672_),
    .C1(_1673_),
    .D1(_1674_),
    .Y(_1675_)
  );
  sky130_fd_sc_hd__or3_2 _4019_ (
    .A(_1647_),
    .B(_1611_),
    .C(_1357_),
    .X(_1676_)
  );
  sky130_fd_sc_hd__or3_2 _4020_ (
    .A(_1649_),
    .B(_1613_),
    .C(_1492_),
    .X(_1677_)
  );
  sky130_fd_sc_hd__or3_2 _4021_ (
    .A(_1651_),
    .B(_1494_),
    .C(_1615_),
    .X(_1678_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4022_ (
    .A1(_1646_),
    .A2(_1610_),
    .B1(_1676_),
    .C1(_1677_),
    .D1(_1678_),
    .Y(_1679_)
  );
  sky130_fd_sc_hd__or4_2 _4023_ (
    .A(_1669_),
    .B(_1671_),
    .C(_1675_),
    .D(_1679_),
    .X(_1680_)
  );
  sky130_fd_sc_hd__or4_2 _4024_ (
    .A(_1657_),
    .B(_1659_),
    .C(_1664_),
    .D(_1680_),
    .X(_1681_)
  );
  sky130_fd_sc_hd__buf_1 _4025_ (
    .A(_1681_),
    .X(\g_bit[20].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _4026_ (
    .A1(\g_bit[21].g_word[30].r_bit.Q ),
    .A2(_1501_),
    .A3(_1502_),
    .B1(_1503_),
    .B2(\g_bit[21].g_word[28].r_bit.Q ),
    .X(_1682_)
  );
  sky130_fd_sc_hd__a221o_2 _4027_ (
    .A1(\g_bit[21].g_word[4].r_bit.Q ),
    .A2(_1499_),
    .B1(_1500_),
    .B2(\g_bit[21].g_word[26].r_bit.Q ),
    .C1(_1682_),
    .X(_1683_)
  );
  sky130_fd_sc_hd__a22o_2 _4028_ (
    .A1(\g_bit[21].g_word[5].r_bit.Q ),
    .A2(_1508_),
    .B1(_1509_),
    .B2(\g_bit[21].g_word[2].r_bit.Q ),
    .X(_1684_)
  );
  sky130_fd_sc_hd__a221o_2 _4029_ (
    .A1(\g_bit[21].g_word[25].r_bit.Q ),
    .A2(_1506_),
    .B1(_1507_),
    .B2(\g_bit[21].g_word[31].r_bit.Q ),
    .C1(_1684_),
    .X(_1685_)
  );
  sky130_fd_sc_hd__a22o_2 _4030_ (
    .A1(\g_bit[21].g_word[13].r_bit.Q ),
    .A2(_1512_),
    .B1(_1513_),
    .B2(\g_bit[21].g_word[15].r_bit.Q ),
    .X(_1686_)
  );
  sky130_fd_sc_hd__a22o_2 _4031_ (
    .A1(\g_bit[21].g_word[11].r_bit.Q ),
    .A2(_1515_),
    .B1(_1516_),
    .B2(\g_bit[21].g_word[20].r_bit.Q ),
    .X(_1687_)
  );
  sky130_fd_sc_hd__a22o_2 _4032_ (
    .A1(\g_bit[21].g_word[19].r_bit.Q ),
    .A2(_1518_),
    .B1(_1519_),
    .B2(\g_bit[21].g_word[21].r_bit.Q ),
    .X(_1688_)
  );
  sky130_fd_sc_hd__a22o_2 _4033_ (
    .A1(\g_bit[21].g_word[17].r_bit.Q ),
    .A2(_1521_),
    .B1(_1522_),
    .B2(\g_bit[21].g_word[12].r_bit.Q ),
    .X(_1689_)
  );
  sky130_fd_sc_hd__or4_2 _4034_ (
    .A(_1686_),
    .B(_1687_),
    .C(_1688_),
    .D(_1689_),
    .X(_1690_)
  );
  sky130_fd_sc_hd__inv_2 _4035_ (
    .A(\g_bit[21].g_word[7].r_bit.Q ),
    .Y(_1691_)
  );
  sky130_fd_sc_hd__nor3_2 _4036_ (
    .A(_1691_),
    .B(_1374_),
    .C(_1440_),
    .Y(_1692_)
  );
  sky130_fd_sc_hd__inv_2 _4037_ (
    .A(\g_bit[21].g_word[3].r_bit.Q ),
    .Y(_1693_)
  );
  sky130_fd_sc_hd__nor3_2 _4038_ (
    .A(_1693_),
    .B(_1529_),
    .C(_1530_),
    .Y(_1694_)
  );
  sky130_fd_sc_hd__and3_2 _4039_ (
    .A(\g_bit[21].g_word[24].r_bit.Q ),
    .B(_1444_),
    .C(_1633_),
    .X(_1695_)
  );
  sky130_fd_sc_hd__a2111o_2 _4040_ (
    .A1(\g_bit[21].g_word[29].r_bit.Q ),
    .A2(_1525_),
    .B1(_1692_),
    .C1(_1694_),
    .D1(_1695_),
    .X(_1696_)
  );
  sky130_fd_sc_hd__and3_2 _4041_ (
    .A(\g_bit[21].g_word[27].r_bit.Q ),
    .B(_1536_),
    .C(_1537_),
    .X(_1697_)
  );
  sky130_fd_sc_hd__a221o_2 _4042_ (
    .A1(\g_bit[21].g_word[6].r_bit.Q ),
    .A2(_1534_),
    .B1(_1535_),
    .B2(\g_bit[21].g_word[1].r_bit.Q ),
    .C1(_1697_),
    .X(_1698_)
  );
  sky130_fd_sc_hd__inv_2 _4043_ (
    .A(\g_bit[21].g_word[23].r_bit.Q ),
    .Y(_1699_)
  );
  sky130_fd_sc_hd__inv_2 _4044_ (
    .A(\g_bit[21].g_word[10].r_bit.Q ),
    .Y(_1700_)
  );
  sky130_fd_sc_hd__or3_2 _4045_ (
    .A(_1700_),
    .B(_1137_),
    .C(_1384_),
    .X(_1701_)
  );
  sky130_fd_sc_hd__inv_2 _4046_ (
    .A(\g_bit[21].g_word[9].r_bit.Q ),
    .Y(_1702_)
  );
  sky130_fd_sc_hd__or3_2 _4047_ (
    .A(_1702_),
    .B(_1261_),
    .C(_1545_),
    .X(_1703_)
  );
  sky130_fd_sc_hd__inv_2 _4048_ (
    .A(\g_bit[21].g_word[8].r_bit.Q ),
    .Y(_1704_)
  );
  sky130_fd_sc_hd__or3_2 _4049_ (
    .A(_1704_),
    .B(_1389_),
    .C(_1548_),
    .X(_1705_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4050_ (
    .A1(_1699_),
    .A2(_1541_),
    .B1(_1701_),
    .C1(_1703_),
    .D1(_1705_),
    .Y(_1706_)
  );
  sky130_fd_sc_hd__inv_2 _4051_ (
    .A(\g_bit[21].g_word[22].r_bit.Q ),
    .Y(_1707_)
  );
  sky130_fd_sc_hd__inv_2 _4052_ (
    .A(\g_bit[21].g_word[16].r_bit.Q ),
    .Y(_1708_)
  );
  sky130_fd_sc_hd__or3_2 _4053_ (
    .A(_1708_),
    .B(_1268_),
    .C(_1554_),
    .X(_1709_)
  );
  sky130_fd_sc_hd__inv_2 _4054_ (
    .A(\g_bit[21].g_word[14].r_bit.Q ),
    .Y(_1710_)
  );
  sky130_fd_sc_hd__or3_2 _4055_ (
    .A(_1710_),
    .B(_1557_),
    .C(_1461_),
    .X(_1711_)
  );
  sky130_fd_sc_hd__inv_2 _4056_ (
    .A(\g_bit[21].g_word[18].r_bit.Q ),
    .Y(_1712_)
  );
  sky130_fd_sc_hd__or3_2 _4057_ (
    .A(_1712_),
    .B(_1464_),
    .C(_1560_),
    .X(_1713_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4058_ (
    .A1(_1707_),
    .A2(_1552_),
    .B1(_1709_),
    .C1(_1711_),
    .D1(_1713_),
    .Y(_1714_)
  );
  sky130_fd_sc_hd__or4_2 _4059_ (
    .A(_1696_),
    .B(_1698_),
    .C(_1706_),
    .D(_1714_),
    .X(_1715_)
  );
  sky130_fd_sc_hd__or4_2 _4060_ (
    .A(_1683_),
    .B(_1685_),
    .C(_1690_),
    .D(_1715_),
    .X(_1716_)
  );
  sky130_fd_sc_hd__buf_1 _4061_ (
    .A(_1716_),
    .X(\g_bit[21].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _4062_ (
    .A1(\g_bit[21].g_word[30].r_bit.Q ),
    .A2(_1567_),
    .A3(_1568_),
    .B1(_1569_),
    .B2(\g_bit[21].g_word[28].r_bit.Q ),
    .X(_1717_)
  );
  sky130_fd_sc_hd__a221o_2 _4063_ (
    .A1(\g_bit[21].g_word[4].r_bit.Q ),
    .A2(_1565_),
    .B1(_1566_),
    .B2(\g_bit[21].g_word[26].r_bit.Q ),
    .C1(_1717_),
    .X(_1718_)
  );
  sky130_fd_sc_hd__a22o_2 _4064_ (
    .A1(\g_bit[21].g_word[5].r_bit.Q ),
    .A2(_1574_),
    .B1(_1575_),
    .B2(\g_bit[21].g_word[2].r_bit.Q ),
    .X(_1719_)
  );
  sky130_fd_sc_hd__a221o_2 _4065_ (
    .A1(\g_bit[21].g_word[25].r_bit.Q ),
    .A2(_1572_),
    .B1(_1573_),
    .B2(\g_bit[21].g_word[31].r_bit.Q ),
    .C1(_1719_),
    .X(_1720_)
  );
  sky130_fd_sc_hd__a22o_2 _4066_ (
    .A1(\g_bit[21].g_word[13].r_bit.Q ),
    .A2(_1578_),
    .B1(_1579_),
    .B2(\g_bit[21].g_word[15].r_bit.Q ),
    .X(_1721_)
  );
  sky130_fd_sc_hd__a22o_2 _4067_ (
    .A1(\g_bit[21].g_word[20].r_bit.Q ),
    .A2(_1581_),
    .B1(_1582_),
    .B2(\g_bit[21].g_word[11].r_bit.Q ),
    .X(_1722_)
  );
  sky130_fd_sc_hd__a22o_2 _4068_ (
    .A1(\g_bit[21].g_word[19].r_bit.Q ),
    .A2(_1584_),
    .B1(_1585_),
    .B2(\g_bit[21].g_word[21].r_bit.Q ),
    .X(_1723_)
  );
  sky130_fd_sc_hd__a22o_2 _4069_ (
    .A1(\g_bit[21].g_word[17].r_bit.Q ),
    .A2(_1587_),
    .B1(_1588_),
    .B2(\g_bit[21].g_word[12].r_bit.Q ),
    .X(_1724_)
  );
  sky130_fd_sc_hd__or4_2 _4070_ (
    .A(_1721_),
    .B(_1722_),
    .C(_1723_),
    .D(_1724_),
    .X(_1725_)
  );
  sky130_fd_sc_hd__nor3_2 _4071_ (
    .A(_1691_),
    .B(_1478_),
    .C(_1411_),
    .Y(_1726_)
  );
  sky130_fd_sc_hd__nor3_2 _4072_ (
    .A(_1693_),
    .B(_1593_),
    .C(_1480_),
    .Y(_1727_)
  );
  sky130_fd_sc_hd__and3_2 _4073_ (
    .A(\g_bit[21].g_word[24].r_bit.Q ),
    .B(_1667_),
    .C(_1482_),
    .X(_1728_)
  );
  sky130_fd_sc_hd__a2111o_2 _4074_ (
    .A1(\g_bit[21].g_word[29].r_bit.Q ),
    .A2(_1591_),
    .B1(_1726_),
    .C1(_1727_),
    .D1(_1728_),
    .X(_1729_)
  );
  sky130_fd_sc_hd__and3_2 _4075_ (
    .A(\g_bit[21].g_word[27].r_bit.Q ),
    .B(_1599_),
    .C(_1600_),
    .X(_1730_)
  );
  sky130_fd_sc_hd__a221o_2 _4076_ (
    .A1(\g_bit[21].g_word[6].r_bit.Q ),
    .A2(_1597_),
    .B1(_1598_),
    .B2(\g_bit[21].g_word[1].r_bit.Q ),
    .C1(_1730_),
    .X(_1731_)
  );
  sky130_fd_sc_hd__or3_2 _4077_ (
    .A(_1700_),
    .B(_1169_),
    .C(_1418_),
    .X(_1732_)
  );
  sky130_fd_sc_hd__or3_2 _4078_ (
    .A(_1702_),
    .B(_1293_),
    .C(_1605_),
    .X(_1733_)
  );
  sky130_fd_sc_hd__or3_2 _4079_ (
    .A(_1704_),
    .B(_1421_),
    .C(_1607_),
    .X(_1734_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4080_ (
    .A1(_1699_),
    .A2(_1603_),
    .B1(_1732_),
    .C1(_1733_),
    .D1(_1734_),
    .Y(_1735_)
  );
  sky130_fd_sc_hd__or3_2 _4081_ (
    .A(_1708_),
    .B(_1611_),
    .C(_1357_),
    .X(_1736_)
  );
  sky130_fd_sc_hd__or3_2 _4082_ (
    .A(_1710_),
    .B(_1613_),
    .C(_1492_),
    .X(_1737_)
  );
  sky130_fd_sc_hd__or3_2 _4083_ (
    .A(_1712_),
    .B(_1494_),
    .C(_1615_),
    .X(_1738_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4084_ (
    .A1(_1707_),
    .A2(_1610_),
    .B1(_1736_),
    .C1(_1737_),
    .D1(_1738_),
    .Y(_1739_)
  );
  sky130_fd_sc_hd__or4_2 _4085_ (
    .A(_1729_),
    .B(_1731_),
    .C(_1735_),
    .D(_1739_),
    .X(_1740_)
  );
  sky130_fd_sc_hd__or4_2 _4086_ (
    .A(_1718_),
    .B(_1720_),
    .C(_1725_),
    .D(_1740_),
    .X(_1741_)
  );
  sky130_fd_sc_hd__buf_1 _4087_ (
    .A(_1741_),
    .X(\g_bit[21].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _4088_ (
    .A1(\g_bit[22].g_word[30].r_bit.Q ),
    .A2(_1501_),
    .A3(_1502_),
    .B1(_1503_),
    .B2(\g_bit[22].g_word[28].r_bit.Q ),
    .X(_1742_)
  );
  sky130_fd_sc_hd__a221o_2 _4089_ (
    .A1(\g_bit[22].g_word[4].r_bit.Q ),
    .A2(_1499_),
    .B1(_1500_),
    .B2(\g_bit[22].g_word[26].r_bit.Q ),
    .C1(_1742_),
    .X(_1743_)
  );
  sky130_fd_sc_hd__a22o_2 _4090_ (
    .A1(\g_bit[22].g_word[5].r_bit.Q ),
    .A2(_1508_),
    .B1(_1509_),
    .B2(\g_bit[22].g_word[2].r_bit.Q ),
    .X(_1744_)
  );
  sky130_fd_sc_hd__a221o_2 _4091_ (
    .A1(\g_bit[22].g_word[25].r_bit.Q ),
    .A2(_1506_),
    .B1(_1507_),
    .B2(\g_bit[22].g_word[31].r_bit.Q ),
    .C1(_1744_),
    .X(_1745_)
  );
  sky130_fd_sc_hd__a22o_2 _4092_ (
    .A1(\g_bit[22].g_word[13].r_bit.Q ),
    .A2(_1512_),
    .B1(_1513_),
    .B2(\g_bit[22].g_word[15].r_bit.Q ),
    .X(_1746_)
  );
  sky130_fd_sc_hd__a22o_2 _4093_ (
    .A1(\g_bit[22].g_word[11].r_bit.Q ),
    .A2(_1515_),
    .B1(_1516_),
    .B2(\g_bit[22].g_word[20].r_bit.Q ),
    .X(_1747_)
  );
  sky130_fd_sc_hd__a22o_2 _4094_ (
    .A1(\g_bit[22].g_word[19].r_bit.Q ),
    .A2(_1518_),
    .B1(_1519_),
    .B2(\g_bit[22].g_word[21].r_bit.Q ),
    .X(_1748_)
  );
  sky130_fd_sc_hd__a22o_2 _4095_ (
    .A1(\g_bit[22].g_word[17].r_bit.Q ),
    .A2(_1521_),
    .B1(_1522_),
    .B2(\g_bit[22].g_word[12].r_bit.Q ),
    .X(_1749_)
  );
  sky130_fd_sc_hd__or4_2 _4096_ (
    .A(_1746_),
    .B(_1747_),
    .C(_1748_),
    .D(_1749_),
    .X(_1750_)
  );
  sky130_fd_sc_hd__inv_2 _4097_ (
    .A(\g_bit[22].g_word[7].r_bit.Q ),
    .Y(_1751_)
  );
  sky130_fd_sc_hd__nor3_2 _4098_ (
    .A(_1751_),
    .B(_1374_),
    .C(_1440_),
    .Y(_1752_)
  );
  sky130_fd_sc_hd__inv_2 _4099_ (
    .A(\g_bit[22].g_word[3].r_bit.Q ),
    .Y(_1753_)
  );
  sky130_fd_sc_hd__nor3_2 _4100_ (
    .A(_1753_),
    .B(_1529_),
    .C(_1530_),
    .Y(_1754_)
  );
  sky130_fd_sc_hd__and3_2 _4101_ (
    .A(\g_bit[22].g_word[24].r_bit.Q ),
    .B(_1444_),
    .C(_1633_),
    .X(_1755_)
  );
  sky130_fd_sc_hd__a2111o_2 _4102_ (
    .A1(\g_bit[22].g_word[29].r_bit.Q ),
    .A2(_1525_),
    .B1(_1752_),
    .C1(_1754_),
    .D1(_1755_),
    .X(_1756_)
  );
  sky130_fd_sc_hd__and3_2 _4103_ (
    .A(\g_bit[22].g_word[27].r_bit.Q ),
    .B(_1536_),
    .C(_1537_),
    .X(_1757_)
  );
  sky130_fd_sc_hd__a221o_2 _4104_ (
    .A1(\g_bit[22].g_word[6].r_bit.Q ),
    .A2(_1534_),
    .B1(_1535_),
    .B2(\g_bit[22].g_word[1].r_bit.Q ),
    .C1(_1757_),
    .X(_1758_)
  );
  sky130_fd_sc_hd__inv_2 _4105_ (
    .A(\g_bit[22].g_word[23].r_bit.Q ),
    .Y(_1759_)
  );
  sky130_fd_sc_hd__inv_2 _4106_ (
    .A(\g_bit[22].g_word[10].r_bit.Q ),
    .Y(_1760_)
  );
  sky130_fd_sc_hd__or3_2 _4107_ (
    .A(_1760_),
    .B(_1137_),
    .C(_1384_),
    .X(_1761_)
  );
  sky130_fd_sc_hd__inv_2 _4108_ (
    .A(\g_bit[22].g_word[9].r_bit.Q ),
    .Y(_1762_)
  );
  sky130_fd_sc_hd__or3_2 _4109_ (
    .A(_1762_),
    .B(_1261_),
    .C(_1545_),
    .X(_1763_)
  );
  sky130_fd_sc_hd__inv_2 _4110_ (
    .A(\g_bit[22].g_word[8].r_bit.Q ),
    .Y(_1764_)
  );
  sky130_fd_sc_hd__or3_2 _4111_ (
    .A(_1764_),
    .B(_1389_),
    .C(_1548_),
    .X(_1765_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4112_ (
    .A1(_1759_),
    .A2(_1541_),
    .B1(_1761_),
    .C1(_1763_),
    .D1(_1765_),
    .Y(_1766_)
  );
  sky130_fd_sc_hd__inv_2 _4113_ (
    .A(\g_bit[22].g_word[22].r_bit.Q ),
    .Y(_1767_)
  );
  sky130_fd_sc_hd__inv_2 _4114_ (
    .A(\g_bit[22].g_word[16].r_bit.Q ),
    .Y(_1768_)
  );
  sky130_fd_sc_hd__or3_2 _4115_ (
    .A(_1768_),
    .B(_1268_),
    .C(_1554_),
    .X(_1769_)
  );
  sky130_fd_sc_hd__inv_2 _4116_ (
    .A(\g_bit[22].g_word[14].r_bit.Q ),
    .Y(_1770_)
  );
  sky130_fd_sc_hd__or3_2 _4117_ (
    .A(_1770_),
    .B(_1557_),
    .C(_1461_),
    .X(_1771_)
  );
  sky130_fd_sc_hd__inv_2 _4118_ (
    .A(\g_bit[22].g_word[18].r_bit.Q ),
    .Y(_1772_)
  );
  sky130_fd_sc_hd__or3_2 _4119_ (
    .A(_1772_),
    .B(_1464_),
    .C(_1560_),
    .X(_1773_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4120_ (
    .A1(_1767_),
    .A2(_1552_),
    .B1(_1769_),
    .C1(_1771_),
    .D1(_1773_),
    .Y(_1774_)
  );
  sky130_fd_sc_hd__or4_2 _4121_ (
    .A(_1756_),
    .B(_1758_),
    .C(_1766_),
    .D(_1774_),
    .X(_1775_)
  );
  sky130_fd_sc_hd__or4_2 _4122_ (
    .A(_1743_),
    .B(_1745_),
    .C(_1750_),
    .D(_1775_),
    .X(_1776_)
  );
  sky130_fd_sc_hd__buf_1 _4123_ (
    .A(_1776_),
    .X(\g_bit[22].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _4124_ (
    .A1(\g_bit[22].g_word[30].r_bit.Q ),
    .A2(_1567_),
    .A3(_1568_),
    .B1(_1569_),
    .B2(\g_bit[22].g_word[28].r_bit.Q ),
    .X(_1777_)
  );
  sky130_fd_sc_hd__a221o_2 _4125_ (
    .A1(\g_bit[22].g_word[4].r_bit.Q ),
    .A2(_1565_),
    .B1(_1566_),
    .B2(\g_bit[22].g_word[26].r_bit.Q ),
    .C1(_1777_),
    .X(_1778_)
  );
  sky130_fd_sc_hd__a22o_2 _4126_ (
    .A1(\g_bit[22].g_word[5].r_bit.Q ),
    .A2(_1574_),
    .B1(_1575_),
    .B2(\g_bit[22].g_word[2].r_bit.Q ),
    .X(_1779_)
  );
  sky130_fd_sc_hd__a221o_2 _4127_ (
    .A1(\g_bit[22].g_word[25].r_bit.Q ),
    .A2(_1572_),
    .B1(_1573_),
    .B2(\g_bit[22].g_word[31].r_bit.Q ),
    .C1(_1779_),
    .X(_1780_)
  );
  sky130_fd_sc_hd__a22o_2 _4128_ (
    .A1(\g_bit[22].g_word[13].r_bit.Q ),
    .A2(_1578_),
    .B1(_1579_),
    .B2(\g_bit[22].g_word[15].r_bit.Q ),
    .X(_1781_)
  );
  sky130_fd_sc_hd__a22o_2 _4129_ (
    .A1(\g_bit[22].g_word[20].r_bit.Q ),
    .A2(_1581_),
    .B1(_1582_),
    .B2(\g_bit[22].g_word[11].r_bit.Q ),
    .X(_1782_)
  );
  sky130_fd_sc_hd__a22o_2 _4130_ (
    .A1(\g_bit[22].g_word[19].r_bit.Q ),
    .A2(_1584_),
    .B1(_1585_),
    .B2(\g_bit[22].g_word[21].r_bit.Q ),
    .X(_1783_)
  );
  sky130_fd_sc_hd__a22o_2 _4131_ (
    .A1(\g_bit[22].g_word[17].r_bit.Q ),
    .A2(_1587_),
    .B1(_1588_),
    .B2(\g_bit[22].g_word[12].r_bit.Q ),
    .X(_1784_)
  );
  sky130_fd_sc_hd__or4_2 _4132_ (
    .A(_1781_),
    .B(_1782_),
    .C(_1783_),
    .D(_1784_),
    .X(_1785_)
  );
  sky130_fd_sc_hd__nor3_2 _4133_ (
    .A(_1751_),
    .B(_1478_),
    .C(_1411_),
    .Y(_1786_)
  );
  sky130_fd_sc_hd__nor3_2 _4134_ (
    .A(_1753_),
    .B(_1593_),
    .C(_1480_),
    .Y(_1787_)
  );
  sky130_fd_sc_hd__and3_2 _4135_ (
    .A(\g_bit[22].g_word[24].r_bit.Q ),
    .B(_1667_),
    .C(_1482_),
    .X(_1788_)
  );
  sky130_fd_sc_hd__a2111o_2 _4136_ (
    .A1(\g_bit[22].g_word[29].r_bit.Q ),
    .A2(_1591_),
    .B1(_1786_),
    .C1(_1787_),
    .D1(_1788_),
    .X(_1789_)
  );
  sky130_fd_sc_hd__and3_2 _4137_ (
    .A(\g_bit[22].g_word[27].r_bit.Q ),
    .B(_1599_),
    .C(_1600_),
    .X(_1790_)
  );
  sky130_fd_sc_hd__a221o_2 _4138_ (
    .A1(\g_bit[22].g_word[6].r_bit.Q ),
    .A2(_1597_),
    .B1(_1598_),
    .B2(\g_bit[22].g_word[1].r_bit.Q ),
    .C1(_1790_),
    .X(_1791_)
  );
  sky130_fd_sc_hd__or3_2 _4139_ (
    .A(_1760_),
    .B(_1169_),
    .C(_1418_),
    .X(_1792_)
  );
  sky130_fd_sc_hd__or3_2 _4140_ (
    .A(_1762_),
    .B(_1293_),
    .C(_1605_),
    .X(_1793_)
  );
  sky130_fd_sc_hd__or3_2 _4141_ (
    .A(_1764_),
    .B(_1421_),
    .C(_1607_),
    .X(_1794_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4142_ (
    .A1(_1759_),
    .A2(_1603_),
    .B1(_1792_),
    .C1(_1793_),
    .D1(_1794_),
    .Y(_1795_)
  );
  sky130_fd_sc_hd__or3_2 _4143_ (
    .A(_1768_),
    .B(_1611_),
    .C(_1357_),
    .X(_1796_)
  );
  sky130_fd_sc_hd__or3_2 _4144_ (
    .A(_1770_),
    .B(_1613_),
    .C(_1492_),
    .X(_1797_)
  );
  sky130_fd_sc_hd__or3_2 _4145_ (
    .A(_1772_),
    .B(_1494_),
    .C(_1615_),
    .X(_1798_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4146_ (
    .A1(_1767_),
    .A2(_1610_),
    .B1(_1796_),
    .C1(_1797_),
    .D1(_1798_),
    .Y(_1799_)
  );
  sky130_fd_sc_hd__or4_2 _4147_ (
    .A(_1789_),
    .B(_1791_),
    .C(_1795_),
    .D(_1799_),
    .X(_1800_)
  );
  sky130_fd_sc_hd__or4_2 _4148_ (
    .A(_1778_),
    .B(_1780_),
    .C(_1785_),
    .D(_1800_),
    .X(_1801_)
  );
  sky130_fd_sc_hd__buf_1 _4149_ (
    .A(_1801_),
    .X(\g_bit[22].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _4150_ (
    .A1(\g_bit[23].g_word[30].r_bit.Q ),
    .A2(_1501_),
    .A3(_1502_),
    .B1(_1503_),
    .B2(\g_bit[23].g_word[28].r_bit.Q ),
    .X(_1802_)
  );
  sky130_fd_sc_hd__a221o_2 _4151_ (
    .A1(\g_bit[23].g_word[4].r_bit.Q ),
    .A2(_1499_),
    .B1(_1500_),
    .B2(\g_bit[23].g_word[26].r_bit.Q ),
    .C1(_1802_),
    .X(_1803_)
  );
  sky130_fd_sc_hd__a22o_2 _4152_ (
    .A1(\g_bit[23].g_word[5].r_bit.Q ),
    .A2(_1508_),
    .B1(_1509_),
    .B2(\g_bit[23].g_word[2].r_bit.Q ),
    .X(_1804_)
  );
  sky130_fd_sc_hd__a221o_2 _4153_ (
    .A1(\g_bit[23].g_word[25].r_bit.Q ),
    .A2(_1506_),
    .B1(_1507_),
    .B2(\g_bit[23].g_word[31].r_bit.Q ),
    .C1(_1804_),
    .X(_1805_)
  );
  sky130_fd_sc_hd__a22o_2 _4154_ (
    .A1(\g_bit[23].g_word[13].r_bit.Q ),
    .A2(_1512_),
    .B1(_1513_),
    .B2(\g_bit[23].g_word[15].r_bit.Q ),
    .X(_1806_)
  );
  sky130_fd_sc_hd__a22o_2 _4155_ (
    .A1(\g_bit[23].g_word[11].r_bit.Q ),
    .A2(_1515_),
    .B1(_1516_),
    .B2(\g_bit[23].g_word[20].r_bit.Q ),
    .X(_1807_)
  );
  sky130_fd_sc_hd__a22o_2 _4156_ (
    .A1(\g_bit[23].g_word[19].r_bit.Q ),
    .A2(_1518_),
    .B1(_1519_),
    .B2(\g_bit[23].g_word[21].r_bit.Q ),
    .X(_1808_)
  );
  sky130_fd_sc_hd__a22o_2 _4157_ (
    .A1(\g_bit[23].g_word[17].r_bit.Q ),
    .A2(_1521_),
    .B1(_1522_),
    .B2(\g_bit[23].g_word[12].r_bit.Q ),
    .X(_1809_)
  );
  sky130_fd_sc_hd__or4_2 _4158_ (
    .A(_1806_),
    .B(_1807_),
    .C(_1808_),
    .D(_1809_),
    .X(_1810_)
  );
  sky130_fd_sc_hd__inv_2 _4159_ (
    .A(\g_bit[23].g_word[7].r_bit.Q ),
    .Y(_1811_)
  );
  sky130_fd_sc_hd__nor3_2 _4160_ (
    .A(_1811_),
    .B(_1374_),
    .C(_1440_),
    .Y(_1812_)
  );
  sky130_fd_sc_hd__inv_2 _4161_ (
    .A(\g_bit[23].g_word[3].r_bit.Q ),
    .Y(_1813_)
  );
  sky130_fd_sc_hd__nor3_2 _4162_ (
    .A(_1813_),
    .B(_1529_),
    .C(_1530_),
    .Y(_1814_)
  );
  sky130_fd_sc_hd__and3_2 _4163_ (
    .A(\g_bit[23].g_word[24].r_bit.Q ),
    .B(_1444_),
    .C(_1633_),
    .X(_1815_)
  );
  sky130_fd_sc_hd__a2111o_2 _4164_ (
    .A1(\g_bit[23].g_word[29].r_bit.Q ),
    .A2(_1525_),
    .B1(_1812_),
    .C1(_1814_),
    .D1(_1815_),
    .X(_1816_)
  );
  sky130_fd_sc_hd__and3_2 _4165_ (
    .A(\g_bit[23].g_word[27].r_bit.Q ),
    .B(_1536_),
    .C(_1537_),
    .X(_1817_)
  );
  sky130_fd_sc_hd__a221o_2 _4166_ (
    .A1(\g_bit[23].g_word[6].r_bit.Q ),
    .A2(_1534_),
    .B1(_1535_),
    .B2(\g_bit[23].g_word[1].r_bit.Q ),
    .C1(_1817_),
    .X(_1818_)
  );
  sky130_fd_sc_hd__inv_2 _4167_ (
    .A(\g_bit[23].g_word[23].r_bit.Q ),
    .Y(_1819_)
  );
  sky130_fd_sc_hd__inv_2 _4168_ (
    .A(\g_bit[23].g_word[10].r_bit.Q ),
    .Y(_1820_)
  );
  sky130_fd_sc_hd__or3_2 _4169_ (
    .A(_1820_),
    .B(_0016_),
    .C(_1384_),
    .X(_1821_)
  );
  sky130_fd_sc_hd__inv_2 _4170_ (
    .A(\g_bit[23].g_word[9].r_bit.Q ),
    .Y(_1822_)
  );
  sky130_fd_sc_hd__or3_2 _4171_ (
    .A(_1822_),
    .B(_1261_),
    .C(_1545_),
    .X(_1823_)
  );
  sky130_fd_sc_hd__inv_2 _4172_ (
    .A(\g_bit[23].g_word[8].r_bit.Q ),
    .Y(_1824_)
  );
  sky130_fd_sc_hd__or3_2 _4173_ (
    .A(_1824_),
    .B(_1389_),
    .C(_1548_),
    .X(_1825_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4174_ (
    .A1(_1819_),
    .A2(_1541_),
    .B1(_1821_),
    .C1(_1823_),
    .D1(_1825_),
    .Y(_1826_)
  );
  sky130_fd_sc_hd__inv_2 _4175_ (
    .A(\g_bit[23].g_word[22].r_bit.Q ),
    .Y(_1827_)
  );
  sky130_fd_sc_hd__inv_2 _4176_ (
    .A(\g_bit[23].g_word[16].r_bit.Q ),
    .Y(_1828_)
  );
  sky130_fd_sc_hd__or3_2 _4177_ (
    .A(_1828_),
    .B(_1268_),
    .C(_1554_),
    .X(_1829_)
  );
  sky130_fd_sc_hd__inv_2 _4178_ (
    .A(\g_bit[23].g_word[14].r_bit.Q ),
    .Y(_1830_)
  );
  sky130_fd_sc_hd__or3_2 _4179_ (
    .A(_1830_),
    .B(_1557_),
    .C(_1461_),
    .X(_1831_)
  );
  sky130_fd_sc_hd__inv_2 _4180_ (
    .A(\g_bit[23].g_word[18].r_bit.Q ),
    .Y(_1832_)
  );
  sky130_fd_sc_hd__or3_2 _4181_ (
    .A(_1832_),
    .B(_1464_),
    .C(_1560_),
    .X(_1833_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4182_ (
    .A1(_1827_),
    .A2(_1552_),
    .B1(_1829_),
    .C1(_1831_),
    .D1(_1833_),
    .Y(_1834_)
  );
  sky130_fd_sc_hd__or4_2 _4183_ (
    .A(_1816_),
    .B(_1818_),
    .C(_1826_),
    .D(_1834_),
    .X(_1835_)
  );
  sky130_fd_sc_hd__or4_2 _4184_ (
    .A(_1803_),
    .B(_1805_),
    .C(_1810_),
    .D(_1835_),
    .X(_1836_)
  );
  sky130_fd_sc_hd__buf_1 _4185_ (
    .A(_1836_),
    .X(\g_bit[23].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _4186_ (
    .A1(\g_bit[23].g_word[30].r_bit.Q ),
    .A2(_1567_),
    .A3(_1568_),
    .B1(_1569_),
    .B2(\g_bit[23].g_word[28].r_bit.Q ),
    .X(_1837_)
  );
  sky130_fd_sc_hd__a221o_2 _4187_ (
    .A1(\g_bit[23].g_word[4].r_bit.Q ),
    .A2(_1565_),
    .B1(_1566_),
    .B2(\g_bit[23].g_word[26].r_bit.Q ),
    .C1(_1837_),
    .X(_1838_)
  );
  sky130_fd_sc_hd__a22o_2 _4188_ (
    .A1(\g_bit[23].g_word[5].r_bit.Q ),
    .A2(_1574_),
    .B1(_1575_),
    .B2(\g_bit[23].g_word[2].r_bit.Q ),
    .X(_1839_)
  );
  sky130_fd_sc_hd__a221o_2 _4189_ (
    .A1(\g_bit[23].g_word[25].r_bit.Q ),
    .A2(_1572_),
    .B1(_1573_),
    .B2(\g_bit[23].g_word[31].r_bit.Q ),
    .C1(_1839_),
    .X(_1840_)
  );
  sky130_fd_sc_hd__a22o_2 _4190_ (
    .A1(\g_bit[23].g_word[13].r_bit.Q ),
    .A2(_1578_),
    .B1(_1579_),
    .B2(\g_bit[23].g_word[15].r_bit.Q ),
    .X(_1841_)
  );
  sky130_fd_sc_hd__a22o_2 _4191_ (
    .A1(\g_bit[23].g_word[20].r_bit.Q ),
    .A2(_1581_),
    .B1(_1582_),
    .B2(\g_bit[23].g_word[11].r_bit.Q ),
    .X(_1842_)
  );
  sky130_fd_sc_hd__a22o_2 _4192_ (
    .A1(\g_bit[23].g_word[19].r_bit.Q ),
    .A2(_1584_),
    .B1(_1585_),
    .B2(\g_bit[23].g_word[21].r_bit.Q ),
    .X(_1843_)
  );
  sky130_fd_sc_hd__a22o_2 _4193_ (
    .A1(\g_bit[23].g_word[17].r_bit.Q ),
    .A2(_1587_),
    .B1(_1588_),
    .B2(\g_bit[23].g_word[12].r_bit.Q ),
    .X(_1844_)
  );
  sky130_fd_sc_hd__or4_2 _4194_ (
    .A(_1841_),
    .B(_1842_),
    .C(_1843_),
    .D(_1844_),
    .X(_1845_)
  );
  sky130_fd_sc_hd__nor3_2 _4195_ (
    .A(_1811_),
    .B(_1478_),
    .C(_1411_),
    .Y(_1846_)
  );
  sky130_fd_sc_hd__nor3_2 _4196_ (
    .A(_1813_),
    .B(_1593_),
    .C(_1480_),
    .Y(_1847_)
  );
  sky130_fd_sc_hd__and3_2 _4197_ (
    .A(\g_bit[23].g_word[24].r_bit.Q ),
    .B(_1667_),
    .C(_1482_),
    .X(_1848_)
  );
  sky130_fd_sc_hd__a2111o_2 _4198_ (
    .A1(\g_bit[23].g_word[29].r_bit.Q ),
    .A2(_1591_),
    .B1(_1846_),
    .C1(_1847_),
    .D1(_1848_),
    .X(_1849_)
  );
  sky130_fd_sc_hd__and3_2 _4199_ (
    .A(\g_bit[23].g_word[27].r_bit.Q ),
    .B(_1599_),
    .C(_1600_),
    .X(_1850_)
  );
  sky130_fd_sc_hd__a221o_2 _4200_ (
    .A1(\g_bit[23].g_word[6].r_bit.Q ),
    .A2(_1597_),
    .B1(_1598_),
    .B2(\g_bit[23].g_word[1].r_bit.Q ),
    .C1(_1850_),
    .X(_1851_)
  );
  sky130_fd_sc_hd__or3_2 _4201_ (
    .A(_1820_),
    .B(_0145_),
    .C(_1418_),
    .X(_1852_)
  );
  sky130_fd_sc_hd__or3_2 _4202_ (
    .A(_1822_),
    .B(_1293_),
    .C(_1605_),
    .X(_1853_)
  );
  sky130_fd_sc_hd__or3_2 _4203_ (
    .A(_1824_),
    .B(_1421_),
    .C(_1607_),
    .X(_1854_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4204_ (
    .A1(_1819_),
    .A2(_1603_),
    .B1(_1852_),
    .C1(_1853_),
    .D1(_1854_),
    .Y(_1855_)
  );
  sky130_fd_sc_hd__or3_2 _4205_ (
    .A(_1828_),
    .B(_1611_),
    .C(_1357_),
    .X(_1856_)
  );
  sky130_fd_sc_hd__or3_2 _4206_ (
    .A(_1830_),
    .B(_1613_),
    .C(_1492_),
    .X(_1857_)
  );
  sky130_fd_sc_hd__or3_2 _4207_ (
    .A(_1832_),
    .B(_1494_),
    .C(_1615_),
    .X(_1858_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4208_ (
    .A1(_1827_),
    .A2(_1610_),
    .B1(_1856_),
    .C1(_1857_),
    .D1(_1858_),
    .Y(_1859_)
  );
  sky130_fd_sc_hd__or4_2 _4209_ (
    .A(_1849_),
    .B(_1851_),
    .C(_1855_),
    .D(_1859_),
    .X(_1860_)
  );
  sky130_fd_sc_hd__or4_2 _4210_ (
    .A(_1838_),
    .B(_1840_),
    .C(_1845_),
    .D(_1860_),
    .X(_1861_)
  );
  sky130_fd_sc_hd__buf_1 _4211_ (
    .A(_1861_),
    .X(\g_bit[23].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _4212_ (
    .A1(\g_bit[24].g_word[30].r_bit.Q ),
    .A2(_1501_),
    .A3(_1502_),
    .B1(_1503_),
    .B2(\g_bit[24].g_word[28].r_bit.Q ),
    .X(_1862_)
  );
  sky130_fd_sc_hd__a221o_2 _4213_ (
    .A1(\g_bit[24].g_word[4].r_bit.Q ),
    .A2(_1499_),
    .B1(_1500_),
    .B2(\g_bit[24].g_word[26].r_bit.Q ),
    .C1(_1862_),
    .X(_1863_)
  );
  sky130_fd_sc_hd__a22o_2 _4214_ (
    .A1(\g_bit[24].g_word[5].r_bit.Q ),
    .A2(_1508_),
    .B1(_1509_),
    .B2(\g_bit[24].g_word[2].r_bit.Q ),
    .X(_1864_)
  );
  sky130_fd_sc_hd__a221o_2 _4215_ (
    .A1(\g_bit[24].g_word[25].r_bit.Q ),
    .A2(_1506_),
    .B1(_1507_),
    .B2(\g_bit[24].g_word[31].r_bit.Q ),
    .C1(_1864_),
    .X(_1865_)
  );
  sky130_fd_sc_hd__a22o_2 _4216_ (
    .A1(\g_bit[24].g_word[13].r_bit.Q ),
    .A2(_1512_),
    .B1(_1513_),
    .B2(\g_bit[24].g_word[15].r_bit.Q ),
    .X(_1866_)
  );
  sky130_fd_sc_hd__a22o_2 _4217_ (
    .A1(\g_bit[24].g_word[11].r_bit.Q ),
    .A2(_1515_),
    .B1(_1516_),
    .B2(\g_bit[24].g_word[20].r_bit.Q ),
    .X(_1867_)
  );
  sky130_fd_sc_hd__a22o_2 _4218_ (
    .A1(\g_bit[24].g_word[19].r_bit.Q ),
    .A2(_1518_),
    .B1(_1519_),
    .B2(\g_bit[24].g_word[21].r_bit.Q ),
    .X(_1868_)
  );
  sky130_fd_sc_hd__a22o_2 _4219_ (
    .A1(\g_bit[24].g_word[17].r_bit.Q ),
    .A2(_1521_),
    .B1(_1522_),
    .B2(\g_bit[24].g_word[12].r_bit.Q ),
    .X(_1869_)
  );
  sky130_fd_sc_hd__or4_2 _4220_ (
    .A(_1866_),
    .B(_1867_),
    .C(_1868_),
    .D(_1869_),
    .X(_1870_)
  );
  sky130_fd_sc_hd__inv_2 _4221_ (
    .A(\g_bit[24].g_word[7].r_bit.Q ),
    .Y(_1871_)
  );
  sky130_fd_sc_hd__nor3_2 _4222_ (
    .A(_1871_),
    .B(_1374_),
    .C(_1440_),
    .Y(_1872_)
  );
  sky130_fd_sc_hd__inv_2 _4223_ (
    .A(\g_bit[24].g_word[3].r_bit.Q ),
    .Y(_1873_)
  );
  sky130_fd_sc_hd__nor3_2 _4224_ (
    .A(_1873_),
    .B(_1529_),
    .C(_1530_),
    .Y(_1874_)
  );
  sky130_fd_sc_hd__and3_2 _4225_ (
    .A(\g_bit[24].g_word[24].r_bit.Q ),
    .B(_1444_),
    .C(_1633_),
    .X(_1875_)
  );
  sky130_fd_sc_hd__a2111o_2 _4226_ (
    .A1(\g_bit[24].g_word[29].r_bit.Q ),
    .A2(_1525_),
    .B1(_1872_),
    .C1(_1874_),
    .D1(_1875_),
    .X(_1876_)
  );
  sky130_fd_sc_hd__and3_2 _4227_ (
    .A(\g_bit[24].g_word[27].r_bit.Q ),
    .B(_1536_),
    .C(_1537_),
    .X(_1877_)
  );
  sky130_fd_sc_hd__a221o_2 _4228_ (
    .A1(\g_bit[24].g_word[6].r_bit.Q ),
    .A2(_1534_),
    .B1(_1535_),
    .B2(\g_bit[24].g_word[1].r_bit.Q ),
    .C1(_1877_),
    .X(_1878_)
  );
  sky130_fd_sc_hd__inv_2 _4229_ (
    .A(\g_bit[24].g_word[23].r_bit.Q ),
    .Y(_1879_)
  );
  sky130_fd_sc_hd__inv_2 _4230_ (
    .A(\g_bit[24].g_word[10].r_bit.Q ),
    .Y(_1880_)
  );
  sky130_fd_sc_hd__or3_2 _4231_ (
    .A(_1880_),
    .B(_0016_),
    .C(_1384_),
    .X(_1881_)
  );
  sky130_fd_sc_hd__inv_2 _4232_ (
    .A(\g_bit[24].g_word[9].r_bit.Q ),
    .Y(_1882_)
  );
  sky130_fd_sc_hd__or3_2 _4233_ (
    .A(_1882_),
    .B(_1261_),
    .C(_1545_),
    .X(_1883_)
  );
  sky130_fd_sc_hd__inv_2 _4234_ (
    .A(\g_bit[24].g_word[8].r_bit.Q ),
    .Y(_1884_)
  );
  sky130_fd_sc_hd__or3_2 _4235_ (
    .A(_1884_),
    .B(_1389_),
    .C(_1548_),
    .X(_1885_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4236_ (
    .A1(_1879_),
    .A2(_1541_),
    .B1(_1881_),
    .C1(_1883_),
    .D1(_1885_),
    .Y(_1886_)
  );
  sky130_fd_sc_hd__inv_2 _4237_ (
    .A(\g_bit[24].g_word[22].r_bit.Q ),
    .Y(_1887_)
  );
  sky130_fd_sc_hd__inv_2 _4238_ (
    .A(\g_bit[24].g_word[16].r_bit.Q ),
    .Y(_1888_)
  );
  sky130_fd_sc_hd__or3_2 _4239_ (
    .A(_1888_),
    .B(_1268_),
    .C(_1554_),
    .X(_1889_)
  );
  sky130_fd_sc_hd__inv_2 _4240_ (
    .A(\g_bit[24].g_word[14].r_bit.Q ),
    .Y(_1890_)
  );
  sky130_fd_sc_hd__or3_2 _4241_ (
    .A(_1890_),
    .B(_1557_),
    .C(_1461_),
    .X(_1891_)
  );
  sky130_fd_sc_hd__inv_2 _4242_ (
    .A(\g_bit[24].g_word[18].r_bit.Q ),
    .Y(_1892_)
  );
  sky130_fd_sc_hd__or3_2 _4243_ (
    .A(_1892_),
    .B(_1464_),
    .C(_1560_),
    .X(_1893_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4244_ (
    .A1(_1887_),
    .A2(_1552_),
    .B1(_1889_),
    .C1(_1891_),
    .D1(_1893_),
    .Y(_1894_)
  );
  sky130_fd_sc_hd__or4_2 _4245_ (
    .A(_1876_),
    .B(_1878_),
    .C(_1886_),
    .D(_1894_),
    .X(_1895_)
  );
  sky130_fd_sc_hd__or4_2 _4246_ (
    .A(_1863_),
    .B(_1865_),
    .C(_1870_),
    .D(_1895_),
    .X(_1896_)
  );
  sky130_fd_sc_hd__buf_1 _4247_ (
    .A(_1896_),
    .X(\g_bit[24].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _4248_ (
    .A1(\g_bit[24].g_word[30].r_bit.Q ),
    .A2(_1567_),
    .A3(_1568_),
    .B1(_1569_),
    .B2(\g_bit[24].g_word[28].r_bit.Q ),
    .X(_1897_)
  );
  sky130_fd_sc_hd__a221o_2 _4249_ (
    .A1(\g_bit[24].g_word[4].r_bit.Q ),
    .A2(_1565_),
    .B1(_1566_),
    .B2(\g_bit[24].g_word[26].r_bit.Q ),
    .C1(_1897_),
    .X(_1898_)
  );
  sky130_fd_sc_hd__a22o_2 _4250_ (
    .A1(\g_bit[24].g_word[5].r_bit.Q ),
    .A2(_1574_),
    .B1(_1575_),
    .B2(\g_bit[24].g_word[2].r_bit.Q ),
    .X(_1899_)
  );
  sky130_fd_sc_hd__a221o_2 _4251_ (
    .A1(\g_bit[24].g_word[25].r_bit.Q ),
    .A2(_1572_),
    .B1(_1573_),
    .B2(\g_bit[24].g_word[31].r_bit.Q ),
    .C1(_1899_),
    .X(_1900_)
  );
  sky130_fd_sc_hd__a22o_2 _4252_ (
    .A1(\g_bit[24].g_word[13].r_bit.Q ),
    .A2(_1578_),
    .B1(_1579_),
    .B2(\g_bit[24].g_word[15].r_bit.Q ),
    .X(_1901_)
  );
  sky130_fd_sc_hd__a22o_2 _4253_ (
    .A1(\g_bit[24].g_word[20].r_bit.Q ),
    .A2(_1581_),
    .B1(_1582_),
    .B2(\g_bit[24].g_word[11].r_bit.Q ),
    .X(_1902_)
  );
  sky130_fd_sc_hd__a22o_2 _4254_ (
    .A1(\g_bit[24].g_word[19].r_bit.Q ),
    .A2(_1584_),
    .B1(_1585_),
    .B2(\g_bit[24].g_word[21].r_bit.Q ),
    .X(_1903_)
  );
  sky130_fd_sc_hd__a22o_2 _4255_ (
    .A1(\g_bit[24].g_word[17].r_bit.Q ),
    .A2(_1587_),
    .B1(_1588_),
    .B2(\g_bit[24].g_word[12].r_bit.Q ),
    .X(_1904_)
  );
  sky130_fd_sc_hd__or4_2 _4256_ (
    .A(_1901_),
    .B(_1902_),
    .C(_1903_),
    .D(_1904_),
    .X(_1905_)
  );
  sky130_fd_sc_hd__nor3_2 _4257_ (
    .A(_1871_),
    .B(_1478_),
    .C(_1411_),
    .Y(_1906_)
  );
  sky130_fd_sc_hd__nor3_2 _4258_ (
    .A(_1873_),
    .B(_1593_),
    .C(_1480_),
    .Y(_1907_)
  );
  sky130_fd_sc_hd__and3_2 _4259_ (
    .A(\g_bit[24].g_word[24].r_bit.Q ),
    .B(_1667_),
    .C(_1482_),
    .X(_1908_)
  );
  sky130_fd_sc_hd__a2111o_2 _4260_ (
    .A1(\g_bit[24].g_word[29].r_bit.Q ),
    .A2(_1591_),
    .B1(_1906_),
    .C1(_1907_),
    .D1(_1908_),
    .X(_1909_)
  );
  sky130_fd_sc_hd__and3_2 _4261_ (
    .A(\g_bit[24].g_word[27].r_bit.Q ),
    .B(_1599_),
    .C(_1600_),
    .X(_1910_)
  );
  sky130_fd_sc_hd__a221o_2 _4262_ (
    .A1(\g_bit[24].g_word[6].r_bit.Q ),
    .A2(_1597_),
    .B1(_1598_),
    .B2(\g_bit[24].g_word[1].r_bit.Q ),
    .C1(_1910_),
    .X(_1911_)
  );
  sky130_fd_sc_hd__or3_2 _4263_ (
    .A(_1880_),
    .B(_0145_),
    .C(_1418_),
    .X(_1912_)
  );
  sky130_fd_sc_hd__or3_2 _4264_ (
    .A(_1882_),
    .B(_1293_),
    .C(_1605_),
    .X(_1913_)
  );
  sky130_fd_sc_hd__or3_2 _4265_ (
    .A(_1884_),
    .B(_1421_),
    .C(_1607_),
    .X(_1914_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4266_ (
    .A1(_1879_),
    .A2(_1603_),
    .B1(_1912_),
    .C1(_1913_),
    .D1(_1914_),
    .Y(_1915_)
  );
  sky130_fd_sc_hd__or3_2 _4267_ (
    .A(_1888_),
    .B(_1611_),
    .C(_1357_),
    .X(_1916_)
  );
  sky130_fd_sc_hd__or3_2 _4268_ (
    .A(_1890_),
    .B(_1613_),
    .C(_1492_),
    .X(_1917_)
  );
  sky130_fd_sc_hd__or3_2 _4269_ (
    .A(_1892_),
    .B(_1494_),
    .C(_1615_),
    .X(_1918_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4270_ (
    .A1(_1887_),
    .A2(_1610_),
    .B1(_1916_),
    .C1(_1917_),
    .D1(_1918_),
    .Y(_1919_)
  );
  sky130_fd_sc_hd__or4_2 _4271_ (
    .A(_1909_),
    .B(_1911_),
    .C(_1915_),
    .D(_1919_),
    .X(_1920_)
  );
  sky130_fd_sc_hd__or4_2 _4272_ (
    .A(_1898_),
    .B(_1900_),
    .C(_1905_),
    .D(_1920_),
    .X(_1921_)
  );
  sky130_fd_sc_hd__buf_1 _4273_ (
    .A(_1921_),
    .X(\g_bit[24].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _4274_ (
    .A1(\g_bit[25].g_word[30].r_bit.Q ),
    .A2(_1501_),
    .A3(_1502_),
    .B1(_1503_),
    .B2(\g_bit[25].g_word[28].r_bit.Q ),
    .X(_1922_)
  );
  sky130_fd_sc_hd__a221o_2 _4275_ (
    .A1(\g_bit[25].g_word[4].r_bit.Q ),
    .A2(_1499_),
    .B1(_1500_),
    .B2(\g_bit[25].g_word[26].r_bit.Q ),
    .C1(_1922_),
    .X(_1923_)
  );
  sky130_fd_sc_hd__a22o_2 _4276_ (
    .A1(\g_bit[25].g_word[5].r_bit.Q ),
    .A2(_1508_),
    .B1(_1509_),
    .B2(\g_bit[25].g_word[2].r_bit.Q ),
    .X(_1924_)
  );
  sky130_fd_sc_hd__a221o_2 _4277_ (
    .A1(\g_bit[25].g_word[25].r_bit.Q ),
    .A2(_1506_),
    .B1(_1507_),
    .B2(\g_bit[25].g_word[31].r_bit.Q ),
    .C1(_1924_),
    .X(_1925_)
  );
  sky130_fd_sc_hd__a22o_2 _4278_ (
    .A1(\g_bit[25].g_word[13].r_bit.Q ),
    .A2(_1512_),
    .B1(_1513_),
    .B2(\g_bit[25].g_word[15].r_bit.Q ),
    .X(_1926_)
  );
  sky130_fd_sc_hd__a22o_2 _4279_ (
    .A1(\g_bit[25].g_word[11].r_bit.Q ),
    .A2(_1515_),
    .B1(_1516_),
    .B2(\g_bit[25].g_word[20].r_bit.Q ),
    .X(_1927_)
  );
  sky130_fd_sc_hd__a22o_2 _4280_ (
    .A1(\g_bit[25].g_word[19].r_bit.Q ),
    .A2(_1518_),
    .B1(_1519_),
    .B2(\g_bit[25].g_word[21].r_bit.Q ),
    .X(_1928_)
  );
  sky130_fd_sc_hd__a22o_2 _4281_ (
    .A1(\g_bit[25].g_word[17].r_bit.Q ),
    .A2(_1521_),
    .B1(_1522_),
    .B2(\g_bit[25].g_word[12].r_bit.Q ),
    .X(_1929_)
  );
  sky130_fd_sc_hd__or4_2 _4282_ (
    .A(_1926_),
    .B(_1927_),
    .C(_1928_),
    .D(_1929_),
    .X(_1930_)
  );
  sky130_fd_sc_hd__inv_2 _4283_ (
    .A(\g_bit[25].g_word[7].r_bit.Q ),
    .Y(_1931_)
  );
  sky130_fd_sc_hd__nor3_2 _4284_ (
    .A(_1931_),
    .B(_1374_),
    .C(_1440_),
    .Y(_1932_)
  );
  sky130_fd_sc_hd__inv_2 _4285_ (
    .A(\g_bit[25].g_word[3].r_bit.Q ),
    .Y(_1933_)
  );
  sky130_fd_sc_hd__nor3_2 _4286_ (
    .A(_1933_),
    .B(_1529_),
    .C(_1530_),
    .Y(_1934_)
  );
  sky130_fd_sc_hd__and3_2 _4287_ (
    .A(\g_bit[25].g_word[24].r_bit.Q ),
    .B(_1444_),
    .C(_1633_),
    .X(_1935_)
  );
  sky130_fd_sc_hd__a2111o_2 _4288_ (
    .A1(\g_bit[25].g_word[29].r_bit.Q ),
    .A2(_1525_),
    .B1(_1932_),
    .C1(_1934_),
    .D1(_1935_),
    .X(_1936_)
  );
  sky130_fd_sc_hd__and3_2 _4289_ (
    .A(\g_bit[25].g_word[27].r_bit.Q ),
    .B(_1536_),
    .C(_1537_),
    .X(_1937_)
  );
  sky130_fd_sc_hd__a221o_2 _4290_ (
    .A1(\g_bit[25].g_word[6].r_bit.Q ),
    .A2(_1534_),
    .B1(_1535_),
    .B2(\g_bit[25].g_word[1].r_bit.Q ),
    .C1(_1937_),
    .X(_1938_)
  );
  sky130_fd_sc_hd__inv_2 _4291_ (
    .A(\g_bit[25].g_word[23].r_bit.Q ),
    .Y(_1939_)
  );
  sky130_fd_sc_hd__inv_2 _4292_ (
    .A(\g_bit[25].g_word[10].r_bit.Q ),
    .Y(_1940_)
  );
  sky130_fd_sc_hd__or3_2 _4293_ (
    .A(_1940_),
    .B(_0016_),
    .C(_1384_),
    .X(_1941_)
  );
  sky130_fd_sc_hd__inv_2 _4294_ (
    .A(\g_bit[25].g_word[9].r_bit.Q ),
    .Y(_1942_)
  );
  sky130_fd_sc_hd__or3_2 _4295_ (
    .A(_1942_),
    .B(_0103_),
    .C(_1545_),
    .X(_1943_)
  );
  sky130_fd_sc_hd__inv_2 _4296_ (
    .A(\g_bit[25].g_word[8].r_bit.Q ),
    .Y(_1944_)
  );
  sky130_fd_sc_hd__or3_2 _4297_ (
    .A(_1944_),
    .B(_1389_),
    .C(_1548_),
    .X(_1945_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4298_ (
    .A1(_1939_),
    .A2(_1541_),
    .B1(_1941_),
    .C1(_1943_),
    .D1(_1945_),
    .Y(_1946_)
  );
  sky130_fd_sc_hd__inv_2 _4299_ (
    .A(\g_bit[25].g_word[22].r_bit.Q ),
    .Y(_1947_)
  );
  sky130_fd_sc_hd__inv_2 _4300_ (
    .A(\g_bit[25].g_word[16].r_bit.Q ),
    .Y(_1948_)
  );
  sky130_fd_sc_hd__or3_2 _4301_ (
    .A(_1948_),
    .B(_0046_),
    .C(_1554_),
    .X(_1949_)
  );
  sky130_fd_sc_hd__inv_2 _4302_ (
    .A(\g_bit[25].g_word[14].r_bit.Q ),
    .Y(_1950_)
  );
  sky130_fd_sc_hd__or3_2 _4303_ (
    .A(_1950_),
    .B(_1557_),
    .C(_1461_),
    .X(_1951_)
  );
  sky130_fd_sc_hd__inv_2 _4304_ (
    .A(\g_bit[25].g_word[18].r_bit.Q ),
    .Y(_1952_)
  );
  sky130_fd_sc_hd__or3_2 _4305_ (
    .A(_1952_),
    .B(_1464_),
    .C(_1560_),
    .X(_1953_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4306_ (
    .A1(_1947_),
    .A2(_1552_),
    .B1(_1949_),
    .C1(_1951_),
    .D1(_1953_),
    .Y(_1954_)
  );
  sky130_fd_sc_hd__or4_2 _4307_ (
    .A(_1936_),
    .B(_1938_),
    .C(_1946_),
    .D(_1954_),
    .X(_1955_)
  );
  sky130_fd_sc_hd__or4_2 _4308_ (
    .A(_1923_),
    .B(_1925_),
    .C(_1930_),
    .D(_1955_),
    .X(_1956_)
  );
  sky130_fd_sc_hd__buf_1 _4309_ (
    .A(_1956_),
    .X(\g_bit[25].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _4310_ (
    .A1(\g_bit[25].g_word[30].r_bit.Q ),
    .A2(_1567_),
    .A3(_1568_),
    .B1(_1569_),
    .B2(\g_bit[25].g_word[28].r_bit.Q ),
    .X(_1957_)
  );
  sky130_fd_sc_hd__a221o_2 _4311_ (
    .A1(\g_bit[25].g_word[4].r_bit.Q ),
    .A2(_1565_),
    .B1(_1566_),
    .B2(\g_bit[25].g_word[26].r_bit.Q ),
    .C1(_1957_),
    .X(_1958_)
  );
  sky130_fd_sc_hd__a22o_2 _4312_ (
    .A1(\g_bit[25].g_word[5].r_bit.Q ),
    .A2(_1574_),
    .B1(_1575_),
    .B2(\g_bit[25].g_word[2].r_bit.Q ),
    .X(_1959_)
  );
  sky130_fd_sc_hd__a221o_2 _4313_ (
    .A1(\g_bit[25].g_word[25].r_bit.Q ),
    .A2(_1572_),
    .B1(_1573_),
    .B2(\g_bit[25].g_word[31].r_bit.Q ),
    .C1(_1959_),
    .X(_1960_)
  );
  sky130_fd_sc_hd__a22o_2 _4314_ (
    .A1(\g_bit[25].g_word[13].r_bit.Q ),
    .A2(_1578_),
    .B1(_1579_),
    .B2(\g_bit[25].g_word[15].r_bit.Q ),
    .X(_1961_)
  );
  sky130_fd_sc_hd__a22o_2 _4315_ (
    .A1(\g_bit[25].g_word[20].r_bit.Q ),
    .A2(_1581_),
    .B1(_1582_),
    .B2(\g_bit[25].g_word[11].r_bit.Q ),
    .X(_1962_)
  );
  sky130_fd_sc_hd__a22o_2 _4316_ (
    .A1(\g_bit[25].g_word[19].r_bit.Q ),
    .A2(_1584_),
    .B1(_1585_),
    .B2(\g_bit[25].g_word[21].r_bit.Q ),
    .X(_1963_)
  );
  sky130_fd_sc_hd__a22o_2 _4317_ (
    .A1(\g_bit[25].g_word[17].r_bit.Q ),
    .A2(_1587_),
    .B1(_1588_),
    .B2(\g_bit[25].g_word[12].r_bit.Q ),
    .X(_1964_)
  );
  sky130_fd_sc_hd__or4_2 _4318_ (
    .A(_1961_),
    .B(_1962_),
    .C(_1963_),
    .D(_1964_),
    .X(_1965_)
  );
  sky130_fd_sc_hd__nor3_2 _4319_ (
    .A(_1931_),
    .B(_1478_),
    .C(_1411_),
    .Y(_1966_)
  );
  sky130_fd_sc_hd__nor3_2 _4320_ (
    .A(_1933_),
    .B(_1593_),
    .C(_1480_),
    .Y(_1967_)
  );
  sky130_fd_sc_hd__and3_2 _4321_ (
    .A(\g_bit[25].g_word[24].r_bit.Q ),
    .B(_1667_),
    .C(_1482_),
    .X(_1968_)
  );
  sky130_fd_sc_hd__a2111o_2 _4322_ (
    .A1(\g_bit[25].g_word[29].r_bit.Q ),
    .A2(_1591_),
    .B1(_1966_),
    .C1(_1967_),
    .D1(_1968_),
    .X(_1969_)
  );
  sky130_fd_sc_hd__and3_2 _4323_ (
    .A(\g_bit[25].g_word[27].r_bit.Q ),
    .B(_1599_),
    .C(_1600_),
    .X(_1970_)
  );
  sky130_fd_sc_hd__a221o_2 _4324_ (
    .A1(\g_bit[25].g_word[6].r_bit.Q ),
    .A2(_1597_),
    .B1(_1598_),
    .B2(\g_bit[25].g_word[1].r_bit.Q ),
    .C1(_1970_),
    .X(_1971_)
  );
  sky130_fd_sc_hd__or3_2 _4325_ (
    .A(_1940_),
    .B(_0145_),
    .C(_1418_),
    .X(_1972_)
  );
  sky130_fd_sc_hd__or3_2 _4326_ (
    .A(_1942_),
    .B(_0227_),
    .C(_1605_),
    .X(_1973_)
  );
  sky130_fd_sc_hd__or3_2 _4327_ (
    .A(_1944_),
    .B(_1421_),
    .C(_1607_),
    .X(_1974_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4328_ (
    .A1(_1939_),
    .A2(_1603_),
    .B1(_1972_),
    .C1(_1973_),
    .D1(_1974_),
    .Y(_1975_)
  );
  sky130_fd_sc_hd__or3_2 _4329_ (
    .A(_1948_),
    .B(_1611_),
    .C(_1357_),
    .X(_1976_)
  );
  sky130_fd_sc_hd__or3_2 _4330_ (
    .A(_1950_),
    .B(_1613_),
    .C(_1492_),
    .X(_1977_)
  );
  sky130_fd_sc_hd__or3_2 _4331_ (
    .A(_1952_),
    .B(_1494_),
    .C(_1615_),
    .X(_1978_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4332_ (
    .A1(_1947_),
    .A2(_1610_),
    .B1(_1976_),
    .C1(_1977_),
    .D1(_1978_),
    .Y(_1979_)
  );
  sky130_fd_sc_hd__or4_2 _4333_ (
    .A(_1969_),
    .B(_1971_),
    .C(_1975_),
    .D(_1979_),
    .X(_1980_)
  );
  sky130_fd_sc_hd__or4_2 _4334_ (
    .A(_1958_),
    .B(_1960_),
    .C(_1965_),
    .D(_1980_),
    .X(_1981_)
  );
  sky130_fd_sc_hd__buf_1 _4335_ (
    .A(_1981_),
    .X(\g_bit[25].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _4336_ (
    .A1(\g_bit[26].g_word[30].r_bit.Q ),
    .A2(_1501_),
    .A3(_1502_),
    .B1(_1503_),
    .B2(\g_bit[26].g_word[28].r_bit.Q ),
    .X(_1982_)
  );
  sky130_fd_sc_hd__a221o_2 _4337_ (
    .A1(\g_bit[26].g_word[4].r_bit.Q ),
    .A2(_1499_),
    .B1(_1500_),
    .B2(\g_bit[26].g_word[26].r_bit.Q ),
    .C1(_1982_),
    .X(_1983_)
  );
  sky130_fd_sc_hd__a22o_2 _4338_ (
    .A1(\g_bit[26].g_word[5].r_bit.Q ),
    .A2(_1508_),
    .B1(_1509_),
    .B2(\g_bit[26].g_word[2].r_bit.Q ),
    .X(_1984_)
  );
  sky130_fd_sc_hd__a221o_2 _4339_ (
    .A1(\g_bit[26].g_word[25].r_bit.Q ),
    .A2(_1506_),
    .B1(_1507_),
    .B2(\g_bit[26].g_word[31].r_bit.Q ),
    .C1(_1984_),
    .X(_1985_)
  );
  sky130_fd_sc_hd__a22o_2 _4340_ (
    .A1(\g_bit[26].g_word[13].r_bit.Q ),
    .A2(_1512_),
    .B1(_1513_),
    .B2(\g_bit[26].g_word[15].r_bit.Q ),
    .X(_1986_)
  );
  sky130_fd_sc_hd__a22o_2 _4341_ (
    .A1(\g_bit[26].g_word[11].r_bit.Q ),
    .A2(_1515_),
    .B1(_1516_),
    .B2(\g_bit[26].g_word[20].r_bit.Q ),
    .X(_1987_)
  );
  sky130_fd_sc_hd__a22o_2 _4342_ (
    .A1(\g_bit[26].g_word[19].r_bit.Q ),
    .A2(_1518_),
    .B1(_1519_),
    .B2(\g_bit[26].g_word[21].r_bit.Q ),
    .X(_1988_)
  );
  sky130_fd_sc_hd__a22o_2 _4343_ (
    .A1(\g_bit[26].g_word[17].r_bit.Q ),
    .A2(_1521_),
    .B1(_1522_),
    .B2(\g_bit[26].g_word[12].r_bit.Q ),
    .X(_1989_)
  );
  sky130_fd_sc_hd__or4_2 _4344_ (
    .A(_1986_),
    .B(_1987_),
    .C(_1988_),
    .D(_1989_),
    .X(_1990_)
  );
  sky130_fd_sc_hd__inv_2 _4345_ (
    .A(\g_bit[26].g_word[7].r_bit.Q ),
    .Y(_1991_)
  );
  sky130_fd_sc_hd__nor3_2 _4346_ (
    .A(_1991_),
    .B(_1374_),
    .C(_1440_),
    .Y(_1992_)
  );
  sky130_fd_sc_hd__inv_2 _4347_ (
    .A(\g_bit[26].g_word[3].r_bit.Q ),
    .Y(_1993_)
  );
  sky130_fd_sc_hd__nor3_2 _4348_ (
    .A(_1993_),
    .B(_1529_),
    .C(_1530_),
    .Y(_1994_)
  );
  sky130_fd_sc_hd__and3_2 _4349_ (
    .A(\g_bit[26].g_word[24].r_bit.Q ),
    .B(_1444_),
    .C(_1633_),
    .X(_1995_)
  );
  sky130_fd_sc_hd__a2111o_2 _4350_ (
    .A1(\g_bit[26].g_word[29].r_bit.Q ),
    .A2(_1525_),
    .B1(_1992_),
    .C1(_1994_),
    .D1(_1995_),
    .X(_1996_)
  );
  sky130_fd_sc_hd__and3_2 _4351_ (
    .A(\g_bit[26].g_word[27].r_bit.Q ),
    .B(_1536_),
    .C(_1537_),
    .X(_1997_)
  );
  sky130_fd_sc_hd__a221o_2 _4352_ (
    .A1(\g_bit[26].g_word[6].r_bit.Q ),
    .A2(_1534_),
    .B1(_1535_),
    .B2(\g_bit[26].g_word[1].r_bit.Q ),
    .C1(_1997_),
    .X(_1998_)
  );
  sky130_fd_sc_hd__inv_2 _4353_ (
    .A(\g_bit[26].g_word[23].r_bit.Q ),
    .Y(_1999_)
  );
  sky130_fd_sc_hd__inv_2 _4354_ (
    .A(\g_bit[26].g_word[10].r_bit.Q ),
    .Y(_2000_)
  );
  sky130_fd_sc_hd__or3_2 _4355_ (
    .A(_2000_),
    .B(_0016_),
    .C(_1384_),
    .X(_2001_)
  );
  sky130_fd_sc_hd__inv_2 _4356_ (
    .A(\g_bit[26].g_word[9].r_bit.Q ),
    .Y(_2002_)
  );
  sky130_fd_sc_hd__or3_2 _4357_ (
    .A(_2002_),
    .B(_0103_),
    .C(_1545_),
    .X(_2003_)
  );
  sky130_fd_sc_hd__inv_2 _4358_ (
    .A(\g_bit[26].g_word[8].r_bit.Q ),
    .Y(_2004_)
  );
  sky130_fd_sc_hd__or3_2 _4359_ (
    .A(_2004_),
    .B(_1389_),
    .C(_1548_),
    .X(_2005_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4360_ (
    .A1(_1999_),
    .A2(_1541_),
    .B1(_2001_),
    .C1(_2003_),
    .D1(_2005_),
    .Y(_2006_)
  );
  sky130_fd_sc_hd__inv_2 _4361_ (
    .A(\g_bit[26].g_word[22].r_bit.Q ),
    .Y(_2007_)
  );
  sky130_fd_sc_hd__inv_2 _4362_ (
    .A(\g_bit[26].g_word[16].r_bit.Q ),
    .Y(_2008_)
  );
  sky130_fd_sc_hd__or3_2 _4363_ (
    .A(_2008_),
    .B(_0046_),
    .C(_1554_),
    .X(_2009_)
  );
  sky130_fd_sc_hd__inv_2 _4364_ (
    .A(\g_bit[26].g_word[14].r_bit.Q ),
    .Y(_2010_)
  );
  sky130_fd_sc_hd__or3_2 _4365_ (
    .A(_2010_),
    .B(_1557_),
    .C(_1461_),
    .X(_2011_)
  );
  sky130_fd_sc_hd__inv_2 _4366_ (
    .A(\g_bit[26].g_word[18].r_bit.Q ),
    .Y(_2012_)
  );
  sky130_fd_sc_hd__or3_2 _4367_ (
    .A(_2012_),
    .B(_1464_),
    .C(_1560_),
    .X(_2013_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4368_ (
    .A1(_2007_),
    .A2(_1552_),
    .B1(_2009_),
    .C1(_2011_),
    .D1(_2013_),
    .Y(_2014_)
  );
  sky130_fd_sc_hd__or4_2 _4369_ (
    .A(_1996_),
    .B(_1998_),
    .C(_2006_),
    .D(_2014_),
    .X(_2015_)
  );
  sky130_fd_sc_hd__or4_2 _4370_ (
    .A(_1983_),
    .B(_1985_),
    .C(_1990_),
    .D(_2015_),
    .X(_2016_)
  );
  sky130_fd_sc_hd__buf_1 _4371_ (
    .A(_2016_),
    .X(\g_bit[26].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _4372_ (
    .A1(\g_bit[26].g_word[30].r_bit.Q ),
    .A2(_1567_),
    .A3(_1568_),
    .B1(_1569_),
    .B2(\g_bit[26].g_word[28].r_bit.Q ),
    .X(_2017_)
  );
  sky130_fd_sc_hd__a221o_2 _4373_ (
    .A1(\g_bit[26].g_word[4].r_bit.Q ),
    .A2(_1565_),
    .B1(_1566_),
    .B2(\g_bit[26].g_word[26].r_bit.Q ),
    .C1(_2017_),
    .X(_2018_)
  );
  sky130_fd_sc_hd__a22o_2 _4374_ (
    .A1(\g_bit[26].g_word[5].r_bit.Q ),
    .A2(_1574_),
    .B1(_1575_),
    .B2(\g_bit[26].g_word[2].r_bit.Q ),
    .X(_2019_)
  );
  sky130_fd_sc_hd__a221o_2 _4375_ (
    .A1(\g_bit[26].g_word[25].r_bit.Q ),
    .A2(_1572_),
    .B1(_1573_),
    .B2(\g_bit[26].g_word[31].r_bit.Q ),
    .C1(_2019_),
    .X(_2020_)
  );
  sky130_fd_sc_hd__a22o_2 _4376_ (
    .A1(\g_bit[26].g_word[13].r_bit.Q ),
    .A2(_1578_),
    .B1(_1579_),
    .B2(\g_bit[26].g_word[15].r_bit.Q ),
    .X(_2021_)
  );
  sky130_fd_sc_hd__a22o_2 _4377_ (
    .A1(\g_bit[26].g_word[20].r_bit.Q ),
    .A2(_1581_),
    .B1(_1582_),
    .B2(\g_bit[26].g_word[11].r_bit.Q ),
    .X(_2022_)
  );
  sky130_fd_sc_hd__a22o_2 _4378_ (
    .A1(\g_bit[26].g_word[19].r_bit.Q ),
    .A2(_1584_),
    .B1(_1585_),
    .B2(\g_bit[26].g_word[21].r_bit.Q ),
    .X(_2023_)
  );
  sky130_fd_sc_hd__a22o_2 _4379_ (
    .A1(\g_bit[26].g_word[17].r_bit.Q ),
    .A2(_1587_),
    .B1(_1588_),
    .B2(\g_bit[26].g_word[12].r_bit.Q ),
    .X(_2024_)
  );
  sky130_fd_sc_hd__or4_2 _4380_ (
    .A(_2021_),
    .B(_2022_),
    .C(_2023_),
    .D(_2024_),
    .X(_2025_)
  );
  sky130_fd_sc_hd__nor3_2 _4381_ (
    .A(_1991_),
    .B(_1478_),
    .C(_1411_),
    .Y(_2026_)
  );
  sky130_fd_sc_hd__nor3_2 _4382_ (
    .A(_1993_),
    .B(_1593_),
    .C(_1480_),
    .Y(_2027_)
  );
  sky130_fd_sc_hd__and3_2 _4383_ (
    .A(\g_bit[26].g_word[24].r_bit.Q ),
    .B(_1667_),
    .C(_1482_),
    .X(_2028_)
  );
  sky130_fd_sc_hd__a2111o_2 _4384_ (
    .A1(\g_bit[26].g_word[29].r_bit.Q ),
    .A2(_1591_),
    .B1(_2026_),
    .C1(_2027_),
    .D1(_2028_),
    .X(_2029_)
  );
  sky130_fd_sc_hd__and3_2 _4385_ (
    .A(\g_bit[26].g_word[27].r_bit.Q ),
    .B(_1599_),
    .C(_1600_),
    .X(_2030_)
  );
  sky130_fd_sc_hd__a221o_2 _4386_ (
    .A1(\g_bit[26].g_word[6].r_bit.Q ),
    .A2(_1597_),
    .B1(_1598_),
    .B2(\g_bit[26].g_word[1].r_bit.Q ),
    .C1(_2030_),
    .X(_2031_)
  );
  sky130_fd_sc_hd__or3_2 _4387_ (
    .A(_2000_),
    .B(_0145_),
    .C(_1418_),
    .X(_2032_)
  );
  sky130_fd_sc_hd__or3_2 _4388_ (
    .A(_2002_),
    .B(_0227_),
    .C(_1605_),
    .X(_2033_)
  );
  sky130_fd_sc_hd__or3_2 _4389_ (
    .A(_2004_),
    .B(_1421_),
    .C(_1607_),
    .X(_2034_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4390_ (
    .A1(_1999_),
    .A2(_1603_),
    .B1(_2032_),
    .C1(_2033_),
    .D1(_2034_),
    .Y(_2035_)
  );
  sky130_fd_sc_hd__or3_2 _4391_ (
    .A(_2008_),
    .B(_1611_),
    .C(_0175_),
    .X(_2036_)
  );
  sky130_fd_sc_hd__or3_2 _4392_ (
    .A(_2010_),
    .B(_1613_),
    .C(_1492_),
    .X(_2037_)
  );
  sky130_fd_sc_hd__or3_2 _4393_ (
    .A(_2012_),
    .B(_1494_),
    .C(_1615_),
    .X(_2038_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4394_ (
    .A1(_2007_),
    .A2(_1610_),
    .B1(_2036_),
    .C1(_2037_),
    .D1(_2038_),
    .Y(_2039_)
  );
  sky130_fd_sc_hd__or4_2 _4395_ (
    .A(_2029_),
    .B(_2031_),
    .C(_2035_),
    .D(_2039_),
    .X(_2040_)
  );
  sky130_fd_sc_hd__or4_2 _4396_ (
    .A(_2018_),
    .B(_2020_),
    .C(_2025_),
    .D(_2040_),
    .X(_2041_)
  );
  sky130_fd_sc_hd__buf_1 _4397_ (
    .A(_2041_),
    .X(\g_bit[26].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _4398_ (
    .A1(\g_bit[27].g_word[30].r_bit.Q ),
    .A2(_1501_),
    .A3(_1502_),
    .B1(_1503_),
    .B2(\g_bit[27].g_word[28].r_bit.Q ),
    .X(_2042_)
  );
  sky130_fd_sc_hd__a221o_2 _4399_ (
    .A1(\g_bit[27].g_word[4].r_bit.Q ),
    .A2(_1499_),
    .B1(_1500_),
    .B2(\g_bit[27].g_word[26].r_bit.Q ),
    .C1(_2042_),
    .X(_2043_)
  );
  sky130_fd_sc_hd__a22o_2 _4400_ (
    .A1(\g_bit[27].g_word[5].r_bit.Q ),
    .A2(_1508_),
    .B1(_1509_),
    .B2(\g_bit[27].g_word[2].r_bit.Q ),
    .X(_2044_)
  );
  sky130_fd_sc_hd__a221o_2 _4401_ (
    .A1(\g_bit[27].g_word[25].r_bit.Q ),
    .A2(_1506_),
    .B1(_1507_),
    .B2(\g_bit[27].g_word[31].r_bit.Q ),
    .C1(_2044_),
    .X(_2045_)
  );
  sky130_fd_sc_hd__a22o_2 _4402_ (
    .A1(\g_bit[27].g_word[13].r_bit.Q ),
    .A2(_1512_),
    .B1(_1513_),
    .B2(\g_bit[27].g_word[15].r_bit.Q ),
    .X(_2046_)
  );
  sky130_fd_sc_hd__a22o_2 _4403_ (
    .A1(\g_bit[27].g_word[11].r_bit.Q ),
    .A2(_1515_),
    .B1(_1516_),
    .B2(\g_bit[27].g_word[20].r_bit.Q ),
    .X(_2047_)
  );
  sky130_fd_sc_hd__a22o_2 _4404_ (
    .A1(\g_bit[27].g_word[19].r_bit.Q ),
    .A2(_1518_),
    .B1(_1519_),
    .B2(\g_bit[27].g_word[21].r_bit.Q ),
    .X(_2048_)
  );
  sky130_fd_sc_hd__a22o_2 _4405_ (
    .A1(\g_bit[27].g_word[17].r_bit.Q ),
    .A2(_1521_),
    .B1(_1522_),
    .B2(\g_bit[27].g_word[12].r_bit.Q ),
    .X(_2049_)
  );
  sky130_fd_sc_hd__or4_2 _4406_ (
    .A(_2046_),
    .B(_2047_),
    .C(_2048_),
    .D(_2049_),
    .X(_2050_)
  );
  sky130_fd_sc_hd__inv_2 _4407_ (
    .A(\g_bit[27].g_word[7].r_bit.Q ),
    .Y(_2051_)
  );
  sky130_fd_sc_hd__nor3_2 _4408_ (
    .A(_2051_),
    .B(_0081_),
    .C(_1440_),
    .Y(_2052_)
  );
  sky130_fd_sc_hd__inv_2 _4409_ (
    .A(\g_bit[27].g_word[3].r_bit.Q ),
    .Y(_2053_)
  );
  sky130_fd_sc_hd__nor3_2 _4410_ (
    .A(_2053_),
    .B(_1529_),
    .C(_1530_),
    .Y(_2054_)
  );
  sky130_fd_sc_hd__and3_2 _4411_ (
    .A(\g_bit[27].g_word[24].r_bit.Q ),
    .B(_1444_),
    .C(_1633_),
    .X(_2055_)
  );
  sky130_fd_sc_hd__a2111o_2 _4412_ (
    .A1(\g_bit[27].g_word[29].r_bit.Q ),
    .A2(_1525_),
    .B1(_2052_),
    .C1(_2054_),
    .D1(_2055_),
    .X(_2056_)
  );
  sky130_fd_sc_hd__and3_2 _4413_ (
    .A(\g_bit[27].g_word[27].r_bit.Q ),
    .B(_1536_),
    .C(_1537_),
    .X(_2057_)
  );
  sky130_fd_sc_hd__a221o_2 _4414_ (
    .A1(\g_bit[27].g_word[6].r_bit.Q ),
    .A2(_1534_),
    .B1(_1535_),
    .B2(\g_bit[27].g_word[1].r_bit.Q ),
    .C1(_2057_),
    .X(_2058_)
  );
  sky130_fd_sc_hd__inv_2 _4415_ (
    .A(\g_bit[27].g_word[23].r_bit.Q ),
    .Y(_2059_)
  );
  sky130_fd_sc_hd__inv_2 _4416_ (
    .A(\g_bit[27].g_word[10].r_bit.Q ),
    .Y(_2060_)
  );
  sky130_fd_sc_hd__or3_2 _4417_ (
    .A(_2060_),
    .B(_0016_),
    .C(_0048_),
    .X(_2061_)
  );
  sky130_fd_sc_hd__inv_2 _4418_ (
    .A(\g_bit[27].g_word[9].r_bit.Q ),
    .Y(_2062_)
  );
  sky130_fd_sc_hd__or3_2 _4419_ (
    .A(_2062_),
    .B(_0103_),
    .C(_1545_),
    .X(_2063_)
  );
  sky130_fd_sc_hd__inv_2 _4420_ (
    .A(\g_bit[27].g_word[8].r_bit.Q ),
    .Y(_2064_)
  );
  sky130_fd_sc_hd__or3_2 _4421_ (
    .A(_2064_),
    .B(_0106_),
    .C(_1548_),
    .X(_2065_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4422_ (
    .A1(_2059_),
    .A2(_1541_),
    .B1(_2061_),
    .C1(_2063_),
    .D1(_2065_),
    .Y(_2066_)
  );
  sky130_fd_sc_hd__inv_2 _4423_ (
    .A(\g_bit[27].g_word[22].r_bit.Q ),
    .Y(_2067_)
  );
  sky130_fd_sc_hd__inv_2 _4424_ (
    .A(\g_bit[27].g_word[16].r_bit.Q ),
    .Y(_2068_)
  );
  sky130_fd_sc_hd__or3_2 _4425_ (
    .A(_2068_),
    .B(_0046_),
    .C(_1554_),
    .X(_2069_)
  );
  sky130_fd_sc_hd__inv_2 _4426_ (
    .A(\g_bit[27].g_word[14].r_bit.Q ),
    .Y(_2070_)
  );
  sky130_fd_sc_hd__or3_2 _4427_ (
    .A(_2070_),
    .B(_1557_),
    .C(_1461_),
    .X(_2071_)
  );
  sky130_fd_sc_hd__inv_2 _4428_ (
    .A(\g_bit[27].g_word[18].r_bit.Q ),
    .Y(_2072_)
  );
  sky130_fd_sc_hd__or3_2 _4429_ (
    .A(_2072_),
    .B(_1464_),
    .C(_1560_),
    .X(_2073_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4430_ (
    .A1(_2067_),
    .A2(_1552_),
    .B1(_2069_),
    .C1(_2071_),
    .D1(_2073_),
    .Y(_2074_)
  );
  sky130_fd_sc_hd__or4_2 _4431_ (
    .A(_2056_),
    .B(_2058_),
    .C(_2066_),
    .D(_2074_),
    .X(_2075_)
  );
  sky130_fd_sc_hd__or4_2 _4432_ (
    .A(_2043_),
    .B(_2045_),
    .C(_2050_),
    .D(_2075_),
    .X(_2076_)
  );
  sky130_fd_sc_hd__buf_1 _4433_ (
    .A(_2076_),
    .X(\g_bit[27].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _4434_ (
    .A1(\g_bit[27].g_word[30].r_bit.Q ),
    .A2(_1567_),
    .A3(_1568_),
    .B1(_1569_),
    .B2(\g_bit[27].g_word[28].r_bit.Q ),
    .X(_2077_)
  );
  sky130_fd_sc_hd__a221o_2 _4435_ (
    .A1(\g_bit[27].g_word[4].r_bit.Q ),
    .A2(_1565_),
    .B1(_1566_),
    .B2(\g_bit[27].g_word[26].r_bit.Q ),
    .C1(_2077_),
    .X(_2078_)
  );
  sky130_fd_sc_hd__a22o_2 _4436_ (
    .A1(\g_bit[27].g_word[5].r_bit.Q ),
    .A2(_1574_),
    .B1(_1575_),
    .B2(\g_bit[27].g_word[2].r_bit.Q ),
    .X(_2079_)
  );
  sky130_fd_sc_hd__a221o_2 _4437_ (
    .A1(\g_bit[27].g_word[25].r_bit.Q ),
    .A2(_1572_),
    .B1(_1573_),
    .B2(\g_bit[27].g_word[31].r_bit.Q ),
    .C1(_2079_),
    .X(_2080_)
  );
  sky130_fd_sc_hd__a22o_2 _4438_ (
    .A1(\g_bit[27].g_word[13].r_bit.Q ),
    .A2(_1578_),
    .B1(_1579_),
    .B2(\g_bit[27].g_word[15].r_bit.Q ),
    .X(_2081_)
  );
  sky130_fd_sc_hd__a22o_2 _4439_ (
    .A1(\g_bit[27].g_word[20].r_bit.Q ),
    .A2(_1581_),
    .B1(_1582_),
    .B2(\g_bit[27].g_word[11].r_bit.Q ),
    .X(_2082_)
  );
  sky130_fd_sc_hd__a22o_2 _4440_ (
    .A1(\g_bit[27].g_word[19].r_bit.Q ),
    .A2(_1584_),
    .B1(_1585_),
    .B2(\g_bit[27].g_word[21].r_bit.Q ),
    .X(_2083_)
  );
  sky130_fd_sc_hd__a22o_2 _4441_ (
    .A1(\g_bit[27].g_word[17].r_bit.Q ),
    .A2(_1587_),
    .B1(_1588_),
    .B2(\g_bit[27].g_word[12].r_bit.Q ),
    .X(_2084_)
  );
  sky130_fd_sc_hd__or4_2 _4442_ (
    .A(_2081_),
    .B(_2082_),
    .C(_2083_),
    .D(_2084_),
    .X(_2085_)
  );
  sky130_fd_sc_hd__nor3_2 _4443_ (
    .A(_2051_),
    .B(_1478_),
    .C(_0209_),
    .Y(_2086_)
  );
  sky130_fd_sc_hd__nor3_2 _4444_ (
    .A(_2053_),
    .B(_1593_),
    .C(_1480_),
    .Y(_2087_)
  );
  sky130_fd_sc_hd__and3_2 _4445_ (
    .A(\g_bit[27].g_word[24].r_bit.Q ),
    .B(_1667_),
    .C(_1482_),
    .X(_2088_)
  );
  sky130_fd_sc_hd__a2111o_2 _4446_ (
    .A1(\g_bit[27].g_word[29].r_bit.Q ),
    .A2(_1591_),
    .B1(_2086_),
    .C1(_2087_),
    .D1(_2088_),
    .X(_2089_)
  );
  sky130_fd_sc_hd__and3_2 _4447_ (
    .A(\g_bit[27].g_word[27].r_bit.Q ),
    .B(_1599_),
    .C(_1600_),
    .X(_2090_)
  );
  sky130_fd_sc_hd__a221o_2 _4448_ (
    .A1(\g_bit[27].g_word[6].r_bit.Q ),
    .A2(_1597_),
    .B1(_1598_),
    .B2(\g_bit[27].g_word[1].r_bit.Q ),
    .C1(_2090_),
    .X(_2091_)
  );
  sky130_fd_sc_hd__or3_2 _4449_ (
    .A(_2060_),
    .B(_0145_),
    .C(_0177_),
    .X(_2092_)
  );
  sky130_fd_sc_hd__or3_2 _4450_ (
    .A(_2062_),
    .B(_0227_),
    .C(_1605_),
    .X(_2093_)
  );
  sky130_fd_sc_hd__or3_2 _4451_ (
    .A(_2064_),
    .B(_0229_),
    .C(_1607_),
    .X(_2094_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4452_ (
    .A1(_2059_),
    .A2(_1603_),
    .B1(_2092_),
    .C1(_2093_),
    .D1(_2094_),
    .Y(_2095_)
  );
  sky130_fd_sc_hd__or3_2 _4453_ (
    .A(_2068_),
    .B(_1611_),
    .C(_0175_),
    .X(_2096_)
  );
  sky130_fd_sc_hd__or3_2 _4454_ (
    .A(_2070_),
    .B(_1613_),
    .C(_1492_),
    .X(_2097_)
  );
  sky130_fd_sc_hd__or3_2 _4455_ (
    .A(_2072_),
    .B(_1494_),
    .C(_1615_),
    .X(_2098_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4456_ (
    .A1(_2067_),
    .A2(_1610_),
    .B1(_2096_),
    .C1(_2097_),
    .D1(_2098_),
    .Y(_2099_)
  );
  sky130_fd_sc_hd__or4_2 _4457_ (
    .A(_2089_),
    .B(_2091_),
    .C(_2095_),
    .D(_2099_),
    .X(_2100_)
  );
  sky130_fd_sc_hd__or4_2 _4458_ (
    .A(_2078_),
    .B(_2080_),
    .C(_2085_),
    .D(_2100_),
    .X(_2101_)
  );
  sky130_fd_sc_hd__buf_1 _4459_ (
    .A(_2101_),
    .X(\g_bit[27].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _4460_ (
    .A1(\g_bit[28].g_word[30].r_bit.Q ),
    .A2(_1501_),
    .A3(_1502_),
    .B1(_1503_),
    .B2(\g_bit[28].g_word[28].r_bit.Q ),
    .X(_2102_)
  );
  sky130_fd_sc_hd__a221o_2 _4461_ (
    .A1(\g_bit[28].g_word[4].r_bit.Q ),
    .A2(_1499_),
    .B1(_1500_),
    .B2(\g_bit[28].g_word[26].r_bit.Q ),
    .C1(_2102_),
    .X(_2103_)
  );
  sky130_fd_sc_hd__a22o_2 _4462_ (
    .A1(\g_bit[28].g_word[5].r_bit.Q ),
    .A2(_1508_),
    .B1(_1509_),
    .B2(\g_bit[28].g_word[2].r_bit.Q ),
    .X(_2104_)
  );
  sky130_fd_sc_hd__a221o_2 _4463_ (
    .A1(\g_bit[28].g_word[25].r_bit.Q ),
    .A2(_1506_),
    .B1(_1507_),
    .B2(\g_bit[28].g_word[31].r_bit.Q ),
    .C1(_2104_),
    .X(_2105_)
  );
  sky130_fd_sc_hd__a22o_2 _4464_ (
    .A1(\g_bit[28].g_word[13].r_bit.Q ),
    .A2(_1512_),
    .B1(_1513_),
    .B2(\g_bit[28].g_word[15].r_bit.Q ),
    .X(_2106_)
  );
  sky130_fd_sc_hd__a22o_2 _4465_ (
    .A1(\g_bit[28].g_word[11].r_bit.Q ),
    .A2(_1515_),
    .B1(_1516_),
    .B2(\g_bit[28].g_word[20].r_bit.Q ),
    .X(_2107_)
  );
  sky130_fd_sc_hd__a22o_2 _4466_ (
    .A1(\g_bit[28].g_word[19].r_bit.Q ),
    .A2(_1518_),
    .B1(_1519_),
    .B2(\g_bit[28].g_word[21].r_bit.Q ),
    .X(_2108_)
  );
  sky130_fd_sc_hd__a22o_2 _4467_ (
    .A1(\g_bit[28].g_word[17].r_bit.Q ),
    .A2(_1521_),
    .B1(_1522_),
    .B2(\g_bit[28].g_word[12].r_bit.Q ),
    .X(_2109_)
  );
  sky130_fd_sc_hd__or4_2 _4468_ (
    .A(_2106_),
    .B(_2107_),
    .C(_2108_),
    .D(_2109_),
    .X(_2110_)
  );
  sky130_fd_sc_hd__inv_2 _4469_ (
    .A(\g_bit[28].g_word[7].r_bit.Q ),
    .Y(_2111_)
  );
  sky130_fd_sc_hd__nor3_2 _4470_ (
    .A(_2111_),
    .B(_0081_),
    .C(_0003_),
    .Y(_2112_)
  );
  sky130_fd_sc_hd__inv_2 _4471_ (
    .A(\g_bit[28].g_word[3].r_bit.Q ),
    .Y(_2113_)
  );
  sky130_fd_sc_hd__nor3_2 _4472_ (
    .A(_2113_),
    .B(_1529_),
    .C(_1530_),
    .Y(_2114_)
  );
  sky130_fd_sc_hd__and3_2 _4473_ (
    .A(\g_bit[28].g_word[24].r_bit.Q ),
    .B(_0077_),
    .C(_1633_),
    .X(_2115_)
  );
  sky130_fd_sc_hd__a2111o_2 _4474_ (
    .A1(\g_bit[28].g_word[29].r_bit.Q ),
    .A2(_1525_),
    .B1(_2112_),
    .C1(_2114_),
    .D1(_2115_),
    .X(_2116_)
  );
  sky130_fd_sc_hd__and3_2 _4475_ (
    .A(\g_bit[28].g_word[27].r_bit.Q ),
    .B(_1536_),
    .C(_1537_),
    .X(_2117_)
  );
  sky130_fd_sc_hd__a221o_2 _4476_ (
    .A1(\g_bit[28].g_word[6].r_bit.Q ),
    .A2(_1534_),
    .B1(_1535_),
    .B2(\g_bit[28].g_word[1].r_bit.Q ),
    .C1(_2117_),
    .X(_2118_)
  );
  sky130_fd_sc_hd__inv_2 _4477_ (
    .A(\g_bit[28].g_word[23].r_bit.Q ),
    .Y(_2119_)
  );
  sky130_fd_sc_hd__inv_2 _4478_ (
    .A(\g_bit[28].g_word[10].r_bit.Q ),
    .Y(_2120_)
  );
  sky130_fd_sc_hd__or3_2 _4479_ (
    .A(_2120_),
    .B(_0016_),
    .C(_0048_),
    .X(_2121_)
  );
  sky130_fd_sc_hd__inv_2 _4480_ (
    .A(\g_bit[28].g_word[9].r_bit.Q ),
    .Y(_2122_)
  );
  sky130_fd_sc_hd__or3_2 _4481_ (
    .A(_2122_),
    .B(_0103_),
    .C(_1545_),
    .X(_2123_)
  );
  sky130_fd_sc_hd__inv_2 _4482_ (
    .A(\g_bit[28].g_word[8].r_bit.Q ),
    .Y(_2124_)
  );
  sky130_fd_sc_hd__or3_2 _4483_ (
    .A(_2124_),
    .B(_0106_),
    .C(_1548_),
    .X(_2125_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4484_ (
    .A1(_2119_),
    .A2(_1541_),
    .B1(_2121_),
    .C1(_2123_),
    .D1(_2125_),
    .Y(_2126_)
  );
  sky130_fd_sc_hd__inv_2 _4485_ (
    .A(\g_bit[28].g_word[22].r_bit.Q ),
    .Y(_2127_)
  );
  sky130_fd_sc_hd__inv_2 _4486_ (
    .A(\g_bit[28].g_word[16].r_bit.Q ),
    .Y(_2128_)
  );
  sky130_fd_sc_hd__or3_2 _4487_ (
    .A(_2128_),
    .B(_0046_),
    .C(_1554_),
    .X(_2129_)
  );
  sky130_fd_sc_hd__inv_2 _4488_ (
    .A(\g_bit[28].g_word[14].r_bit.Q ),
    .Y(_2130_)
  );
  sky130_fd_sc_hd__or3_2 _4489_ (
    .A(_2130_),
    .B(_1557_),
    .C(_0028_),
    .X(_2131_)
  );
  sky130_fd_sc_hd__inv_2 _4490_ (
    .A(\g_bit[28].g_word[18].r_bit.Q ),
    .Y(_2132_)
  );
  sky130_fd_sc_hd__or3_2 _4491_ (
    .A(_2132_),
    .B(_0118_),
    .C(_1560_),
    .X(_2133_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4492_ (
    .A1(_2127_),
    .A2(_1552_),
    .B1(_2129_),
    .C1(_2131_),
    .D1(_2133_),
    .Y(_2134_)
  );
  sky130_fd_sc_hd__or4_2 _4493_ (
    .A(_2116_),
    .B(_2118_),
    .C(_2126_),
    .D(_2134_),
    .X(_2135_)
  );
  sky130_fd_sc_hd__or4_2 _4494_ (
    .A(_2103_),
    .B(_2105_),
    .C(_2110_),
    .D(_2135_),
    .X(_2136_)
  );
  sky130_fd_sc_hd__buf_1 _4495_ (
    .A(_2136_),
    .X(\g_bit[28].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _4496_ (
    .A1(\g_bit[28].g_word[30].r_bit.Q ),
    .A2(_1567_),
    .A3(_1568_),
    .B1(_1569_),
    .B2(\g_bit[28].g_word[28].r_bit.Q ),
    .X(_2137_)
  );
  sky130_fd_sc_hd__a221o_2 _4497_ (
    .A1(\g_bit[28].g_word[4].r_bit.Q ),
    .A2(_1565_),
    .B1(_1566_),
    .B2(\g_bit[28].g_word[26].r_bit.Q ),
    .C1(_2137_),
    .X(_2138_)
  );
  sky130_fd_sc_hd__a22o_2 _4498_ (
    .A1(\g_bit[28].g_word[5].r_bit.Q ),
    .A2(_1574_),
    .B1(_1575_),
    .B2(\g_bit[28].g_word[2].r_bit.Q ),
    .X(_2139_)
  );
  sky130_fd_sc_hd__a221o_2 _4499_ (
    .A1(\g_bit[28].g_word[25].r_bit.Q ),
    .A2(_1572_),
    .B1(_1573_),
    .B2(\g_bit[28].g_word[31].r_bit.Q ),
    .C1(_2139_),
    .X(_2140_)
  );
  sky130_fd_sc_hd__a22o_2 _4500_ (
    .A1(\g_bit[28].g_word[13].r_bit.Q ),
    .A2(_1578_),
    .B1(_1579_),
    .B2(\g_bit[28].g_word[15].r_bit.Q ),
    .X(_2141_)
  );
  sky130_fd_sc_hd__a22o_2 _4501_ (
    .A1(\g_bit[28].g_word[20].r_bit.Q ),
    .A2(_1581_),
    .B1(_1582_),
    .B2(\g_bit[28].g_word[11].r_bit.Q ),
    .X(_2142_)
  );
  sky130_fd_sc_hd__a22o_2 _4502_ (
    .A1(\g_bit[28].g_word[19].r_bit.Q ),
    .A2(_1584_),
    .B1(_1585_),
    .B2(\g_bit[28].g_word[21].r_bit.Q ),
    .X(_2143_)
  );
  sky130_fd_sc_hd__a22o_2 _4503_ (
    .A1(\g_bit[28].g_word[17].r_bit.Q ),
    .A2(_1587_),
    .B1(_1588_),
    .B2(\g_bit[28].g_word[12].r_bit.Q ),
    .X(_2144_)
  );
  sky130_fd_sc_hd__or4_2 _4504_ (
    .A(_2141_),
    .B(_2142_),
    .C(_2143_),
    .D(_2144_),
    .X(_2145_)
  );
  sky130_fd_sc_hd__nor3_2 _4505_ (
    .A(_2111_),
    .B(_0132_),
    .C(_0209_),
    .Y(_2146_)
  );
  sky130_fd_sc_hd__nor3_2 _4506_ (
    .A(_2113_),
    .B(_1593_),
    .C(_0294_),
    .Y(_2147_)
  );
  sky130_fd_sc_hd__and3_2 _4507_ (
    .A(\g_bit[28].g_word[24].r_bit.Q ),
    .B(_1667_),
    .C(_0207_),
    .X(_2148_)
  );
  sky130_fd_sc_hd__a2111o_2 _4508_ (
    .A1(\g_bit[28].g_word[29].r_bit.Q ),
    .A2(_1591_),
    .B1(_2146_),
    .C1(_2147_),
    .D1(_2148_),
    .X(_2149_)
  );
  sky130_fd_sc_hd__and3_2 _4509_ (
    .A(\g_bit[28].g_word[27].r_bit.Q ),
    .B(_1599_),
    .C(_1600_),
    .X(_2150_)
  );
  sky130_fd_sc_hd__a221o_2 _4510_ (
    .A1(\g_bit[28].g_word[6].r_bit.Q ),
    .A2(_1597_),
    .B1(_1598_),
    .B2(\g_bit[28].g_word[1].r_bit.Q ),
    .C1(_2150_),
    .X(_2151_)
  );
  sky130_fd_sc_hd__or3_2 _4511_ (
    .A(_2120_),
    .B(_0145_),
    .C(_0177_),
    .X(_2152_)
  );
  sky130_fd_sc_hd__or3_2 _4512_ (
    .A(_2122_),
    .B(_0227_),
    .C(_1605_),
    .X(_2153_)
  );
  sky130_fd_sc_hd__or3_2 _4513_ (
    .A(_2124_),
    .B(_0229_),
    .C(_1607_),
    .X(_2154_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4514_ (
    .A1(_2119_),
    .A2(_1603_),
    .B1(_2152_),
    .C1(_2153_),
    .D1(_2154_),
    .Y(_2155_)
  );
  sky130_fd_sc_hd__or3_2 _4515_ (
    .A(_2128_),
    .B(_1611_),
    .C(_0175_),
    .X(_2156_)
  );
  sky130_fd_sc_hd__or3_2 _4516_ (
    .A(_2130_),
    .B(_1613_),
    .C(_0157_),
    .X(_2157_)
  );
  sky130_fd_sc_hd__or3_2 _4517_ (
    .A(_2132_),
    .B(_0240_),
    .C(_1615_),
    .X(_2158_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4518_ (
    .A1(_2127_),
    .A2(_1610_),
    .B1(_2156_),
    .C1(_2157_),
    .D1(_2158_),
    .Y(_2159_)
  );
  sky130_fd_sc_hd__or4_2 _4519_ (
    .A(_2149_),
    .B(_2151_),
    .C(_2155_),
    .D(_2159_),
    .X(_2160_)
  );
  sky130_fd_sc_hd__or4_2 _4520_ (
    .A(_2138_),
    .B(_2140_),
    .C(_2145_),
    .D(_2160_),
    .X(_2161_)
  );
  sky130_fd_sc_hd__buf_1 _4521_ (
    .A(_2161_),
    .X(\g_bit[28].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _4522_ (
    .A1(\g_bit[29].g_word[30].r_bit.Q ),
    .A2(_0022_),
    .A3(_0024_),
    .B1(_0029_),
    .B2(\g_bit[29].g_word[28].r_bit.Q ),
    .X(_2162_)
  );
  sky130_fd_sc_hd__a221o_2 _4523_ (
    .A1(\g_bit[29].g_word[4].r_bit.Q ),
    .A2(_0013_),
    .B1(_0020_),
    .B2(\g_bit[29].g_word[26].r_bit.Q ),
    .C1(_2162_),
    .X(_2163_)
  );
  sky130_fd_sc_hd__a22o_2 _4524_ (
    .A1(\g_bit[29].g_word[5].r_bit.Q ),
    .A2(_0042_),
    .B1(_0049_),
    .B2(\g_bit[29].g_word[2].r_bit.Q ),
    .X(_2164_)
  );
  sky130_fd_sc_hd__a221o_2 _4525_ (
    .A1(\g_bit[29].g_word[25].r_bit.Q ),
    .A2(_0034_),
    .B1(_0038_),
    .B2(\g_bit[29].g_word[31].r_bit.Q ),
    .C1(_2164_),
    .X(_2165_)
  );
  sky130_fd_sc_hd__a22o_2 _4526_ (
    .A1(\g_bit[29].g_word[13].r_bit.Q ),
    .A2(_0053_),
    .B1(_0056_),
    .B2(\g_bit[29].g_word[15].r_bit.Q ),
    .X(_2166_)
  );
  sky130_fd_sc_hd__a22o_2 _4527_ (
    .A1(\g_bit[29].g_word[11].r_bit.Q ),
    .A2(_0059_),
    .B1(_0061_),
    .B2(\g_bit[29].g_word[20].r_bit.Q ),
    .X(_2167_)
  );
  sky130_fd_sc_hd__a22o_2 _4528_ (
    .A1(\g_bit[29].g_word[19].r_bit.Q ),
    .A2(_0064_),
    .B1(_0066_),
    .B2(\g_bit[29].g_word[21].r_bit.Q ),
    .X(_2168_)
  );
  sky130_fd_sc_hd__a22o_2 _4529_ (
    .A1(\g_bit[29].g_word[17].r_bit.Q ),
    .A2(_0069_),
    .B1(_0071_),
    .B2(\g_bit[29].g_word[12].r_bit.Q ),
    .X(_2169_)
  );
  sky130_fd_sc_hd__or4_2 _4530_ (
    .A(_2166_),
    .B(_2167_),
    .C(_2168_),
    .D(_2169_),
    .X(_2170_)
  );
  sky130_fd_sc_hd__inv_2 _4531_ (
    .A(\g_bit[29].g_word[7].r_bit.Q ),
    .Y(_2171_)
  );
  sky130_fd_sc_hd__nor3_2 _4532_ (
    .A(_2171_),
    .B(_0081_),
    .C(_0003_),
    .Y(_2172_)
  );
  sky130_fd_sc_hd__inv_2 _4533_ (
    .A(\g_bit[29].g_word[3].r_bit.Q ),
    .Y(_2173_)
  );
  sky130_fd_sc_hd__nor3_2 _4534_ (
    .A(_2173_),
    .B(_0280_),
    .C(_0082_),
    .Y(_2174_)
  );
  sky130_fd_sc_hd__and3_2 _4535_ (
    .A(\g_bit[29].g_word[24].r_bit.Q ),
    .B(_0077_),
    .C(_1633_),
    .X(_2175_)
  );
  sky130_fd_sc_hd__a2111o_2 _4536_ (
    .A1(\g_bit[29].g_word[29].r_bit.Q ),
    .A2(_0075_),
    .B1(_2172_),
    .C1(_2174_),
    .D1(_2175_),
    .X(_2176_)
  );
  sky130_fd_sc_hd__and3_2 _4537_ (
    .A(\g_bit[29].g_word[27].r_bit.Q ),
    .B(_0093_),
    .C(_0260_),
    .X(_2177_)
  );
  sky130_fd_sc_hd__a221o_2 _4538_ (
    .A1(\g_bit[29].g_word[6].r_bit.Q ),
    .A2(_0089_),
    .B1(_0091_),
    .B2(\g_bit[29].g_word[1].r_bit.Q ),
    .C1(_2177_),
    .X(_2178_)
  );
  sky130_fd_sc_hd__inv_2 _4539_ (
    .A(\g_bit[29].g_word[23].r_bit.Q ),
    .Y(_2179_)
  );
  sky130_fd_sc_hd__inv_2 _4540_ (
    .A(\g_bit[29].g_word[10].r_bit.Q ),
    .Y(_2180_)
  );
  sky130_fd_sc_hd__or3_2 _4541_ (
    .A(_2180_),
    .B(_0016_),
    .C(_0048_),
    .X(_2181_)
  );
  sky130_fd_sc_hd__inv_2 _4542_ (
    .A(\g_bit[29].g_word[9].r_bit.Q ),
    .Y(_2182_)
  );
  sky130_fd_sc_hd__or3_2 _4543_ (
    .A(_2182_),
    .B(_0103_),
    .C(_0041_),
    .X(_2183_)
  );
  sky130_fd_sc_hd__inv_2 _4544_ (
    .A(\g_bit[29].g_word[8].r_bit.Q ),
    .Y(_2184_)
  );
  sky130_fd_sc_hd__or3_2 _4545_ (
    .A(_2184_),
    .B(_0106_),
    .C(_0011_),
    .X(_2185_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4546_ (
    .A1(_2179_),
    .A2(_0100_),
    .B1(_2181_),
    .C1(_2183_),
    .D1(_2185_),
    .Y(_2186_)
  );
  sky130_fd_sc_hd__inv_2 _4547_ (
    .A(\g_bit[29].g_word[22].r_bit.Q ),
    .Y(_2187_)
  );
  sky130_fd_sc_hd__inv_2 _4548_ (
    .A(\g_bit[29].g_word[16].r_bit.Q ),
    .Y(_2188_)
  );
  sky130_fd_sc_hd__or3_2 _4549_ (
    .A(_2188_),
    .B(_0046_),
    .C(_0026_),
    .X(_2189_)
  );
  sky130_fd_sc_hd__inv_2 _4550_ (
    .A(\g_bit[29].g_word[14].r_bit.Q ),
    .Y(_2190_)
  );
  sky130_fd_sc_hd__or3_2 _4551_ (
    .A(_2190_),
    .B(_0107_),
    .C(_0028_),
    .X(_2191_)
  );
  sky130_fd_sc_hd__inv_2 _4552_ (
    .A(\g_bit[29].g_word[18].r_bit.Q ),
    .Y(_2192_)
  );
  sky130_fd_sc_hd__or3_2 _4553_ (
    .A(_2192_),
    .B(_0118_),
    .C(_0018_),
    .X(_2193_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4554_ (
    .A1(_2187_),
    .A2(_0115_),
    .B1(_2189_),
    .C1(_2191_),
    .D1(_2193_),
    .Y(_2194_)
  );
  sky130_fd_sc_hd__or4_2 _4555_ (
    .A(_2176_),
    .B(_2178_),
    .C(_2186_),
    .D(_2194_),
    .X(_2195_)
  );
  sky130_fd_sc_hd__or4_2 _4556_ (
    .A(_2163_),
    .B(_2165_),
    .C(_2170_),
    .D(_2195_),
    .X(_2196_)
  );
  sky130_fd_sc_hd__buf_1 _4557_ (
    .A(_2196_),
    .X(\g_bit[29].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _4558_ (
    .A1(\g_bit[29].g_word[30].r_bit.Q ),
    .A2(_0151_),
    .A3(_0153_),
    .B1(_0158_),
    .B2(\g_bit[29].g_word[28].r_bit.Q ),
    .X(_2197_)
  );
  sky130_fd_sc_hd__a221o_2 _4559_ (
    .A1(\g_bit[29].g_word[4].r_bit.Q ),
    .A2(_0142_),
    .B1(_0149_),
    .B2(\g_bit[29].g_word[26].r_bit.Q ),
    .C1(_2197_),
    .X(_2198_)
  );
  sky130_fd_sc_hd__a22o_2 _4560_ (
    .A1(\g_bit[29].g_word[5].r_bit.Q ),
    .A2(_0171_),
    .B1(_0178_),
    .B2(\g_bit[29].g_word[2].r_bit.Q ),
    .X(_2199_)
  );
  sky130_fd_sc_hd__a221o_2 _4561_ (
    .A1(\g_bit[29].g_word[25].r_bit.Q ),
    .A2(_0163_),
    .B1(_0167_),
    .B2(\g_bit[29].g_word[31].r_bit.Q ),
    .C1(_2199_),
    .X(_2200_)
  );
  sky130_fd_sc_hd__a22o_2 _4562_ (
    .A1(\g_bit[29].g_word[13].r_bit.Q ),
    .A2(_0182_),
    .B1(_0185_),
    .B2(\g_bit[29].g_word[15].r_bit.Q ),
    .X(_2201_)
  );
  sky130_fd_sc_hd__a22o_2 _4563_ (
    .A1(\g_bit[29].g_word[20].r_bit.Q ),
    .A2(_0188_),
    .B1(_0190_),
    .B2(\g_bit[29].g_word[11].r_bit.Q ),
    .X(_2202_)
  );
  sky130_fd_sc_hd__a22o_2 _4564_ (
    .A1(\g_bit[29].g_word[19].r_bit.Q ),
    .A2(_0193_),
    .B1(_0195_),
    .B2(\g_bit[29].g_word[21].r_bit.Q ),
    .X(_2203_)
  );
  sky130_fd_sc_hd__a22o_2 _4565_ (
    .A1(\g_bit[29].g_word[17].r_bit.Q ),
    .A2(_0198_),
    .B1(_0200_),
    .B2(\g_bit[29].g_word[12].r_bit.Q ),
    .X(_2204_)
  );
  sky130_fd_sc_hd__or4_2 _4566_ (
    .A(_2201_),
    .B(_2202_),
    .C(_2203_),
    .D(_2204_),
    .X(_2205_)
  );
  sky130_fd_sc_hd__nor3_2 _4567_ (
    .A(_2171_),
    .B(_0132_),
    .C(_0209_),
    .Y(_2206_)
  );
  sky130_fd_sc_hd__nor3_2 _4568_ (
    .A(_2173_),
    .B(_0309_),
    .C(_0294_),
    .Y(_2207_)
  );
  sky130_fd_sc_hd__and3_2 _4569_ (
    .A(\g_bit[29].g_word[24].r_bit.Q ),
    .B(_1667_),
    .C(_0207_),
    .X(_2208_)
  );
  sky130_fd_sc_hd__a2111o_2 _4570_ (
    .A1(\g_bit[29].g_word[29].r_bit.Q ),
    .A2(_0204_),
    .B1(_2206_),
    .C1(_2207_),
    .D1(_2208_),
    .X(_2209_)
  );
  sky130_fd_sc_hd__and3_2 _4571_ (
    .A(\g_bit[29].g_word[27].r_bit.Q ),
    .B(_0219_),
    .C(_0298_),
    .X(_2210_)
  );
  sky130_fd_sc_hd__a221o_2 _4572_ (
    .A1(\g_bit[29].g_word[6].r_bit.Q ),
    .A2(_0215_),
    .B1(_0217_),
    .B2(\g_bit[29].g_word[1].r_bit.Q ),
    .C1(_2210_),
    .X(_2211_)
  );
  sky130_fd_sc_hd__or3_2 _4573_ (
    .A(_2180_),
    .B(_0145_),
    .C(_0177_),
    .X(_2212_)
  );
  sky130_fd_sc_hd__or3_2 _4574_ (
    .A(_2182_),
    .B(_0227_),
    .C(_0170_),
    .X(_2213_)
  );
  sky130_fd_sc_hd__or3_2 _4575_ (
    .A(_2184_),
    .B(_0229_),
    .C(_0140_),
    .X(_2214_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4576_ (
    .A1(_2179_),
    .A2(_0225_),
    .B1(_2212_),
    .C1(_2213_),
    .D1(_2214_),
    .Y(_2215_)
  );
  sky130_fd_sc_hd__or3_2 _4577_ (
    .A(_2188_),
    .B(_0155_),
    .C(_0175_),
    .X(_2216_)
  );
  sky130_fd_sc_hd__or3_2 _4578_ (
    .A(_2190_),
    .B(_0230_),
    .C(_0157_),
    .X(_2217_)
  );
  sky130_fd_sc_hd__or3_2 _4579_ (
    .A(_2192_),
    .B(_0240_),
    .C(_0147_),
    .X(_2218_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4580_ (
    .A1(_2187_),
    .A2(_0236_),
    .B1(_2216_),
    .C1(_2217_),
    .D1(_2218_),
    .Y(_2219_)
  );
  sky130_fd_sc_hd__or4_2 _4581_ (
    .A(_2209_),
    .B(_2211_),
    .C(_2215_),
    .D(_2219_),
    .X(_2220_)
  );
  sky130_fd_sc_hd__or4_2 _4582_ (
    .A(_2198_),
    .B(_2200_),
    .C(_2205_),
    .D(_2220_),
    .X(_2221_)
  );
  sky130_fd_sc_hd__buf_1 _4583_ (
    .A(_2221_),
    .X(\g_bit[29].r_rs2.D )
  );
  sky130_fd_sc_hd__a32o_2 _4584_ (
    .A1(\g_bit[30].g_word[30].r_bit.Q ),
    .A2(_0022_),
    .A3(_0024_),
    .B1(_0029_),
    .B2(\g_bit[30].g_word[28].r_bit.Q ),
    .X(_2222_)
  );
  sky130_fd_sc_hd__a221o_2 _4585_ (
    .A1(\g_bit[30].g_word[4].r_bit.Q ),
    .A2(_0013_),
    .B1(_0020_),
    .B2(\g_bit[30].g_word[26].r_bit.Q ),
    .C1(_2222_),
    .X(_2223_)
  );
  sky130_fd_sc_hd__a22o_2 _4586_ (
    .A1(\g_bit[30].g_word[5].r_bit.Q ),
    .A2(_0042_),
    .B1(_0049_),
    .B2(\g_bit[30].g_word[2].r_bit.Q ),
    .X(_2224_)
  );
  sky130_fd_sc_hd__a221o_2 _4587_ (
    .A1(\g_bit[30].g_word[25].r_bit.Q ),
    .A2(_0034_),
    .B1(_0038_),
    .B2(\g_bit[30].g_word[31].r_bit.Q ),
    .C1(_2224_),
    .X(_2225_)
  );
  sky130_fd_sc_hd__a22o_2 _4588_ (
    .A1(\g_bit[30].g_word[13].r_bit.Q ),
    .A2(_0053_),
    .B1(_0056_),
    .B2(\g_bit[30].g_word[15].r_bit.Q ),
    .X(_2226_)
  );
  sky130_fd_sc_hd__a22o_2 _4589_ (
    .A1(\g_bit[30].g_word[11].r_bit.Q ),
    .A2(_0059_),
    .B1(_0061_),
    .B2(\g_bit[30].g_word[20].r_bit.Q ),
    .X(_2227_)
  );
  sky130_fd_sc_hd__a22o_2 _4590_ (
    .A1(\g_bit[30].g_word[19].r_bit.Q ),
    .A2(_0064_),
    .B1(_0066_),
    .B2(\g_bit[30].g_word[21].r_bit.Q ),
    .X(_2228_)
  );
  sky130_fd_sc_hd__a22o_2 _4591_ (
    .A1(\g_bit[30].g_word[17].r_bit.Q ),
    .A2(_0069_),
    .B1(_0071_),
    .B2(\g_bit[30].g_word[12].r_bit.Q ),
    .X(_2229_)
  );
  sky130_fd_sc_hd__or4_2 _4592_ (
    .A(_2226_),
    .B(_2227_),
    .C(_2228_),
    .D(_2229_),
    .X(_2230_)
  );
  sky130_fd_sc_hd__inv_2 _4593_ (
    .A(\g_bit[30].g_word[7].r_bit.Q ),
    .Y(_2231_)
  );
  sky130_fd_sc_hd__nor3_2 _4594_ (
    .A(_2231_),
    .B(_0081_),
    .C(_0003_),
    .Y(_2232_)
  );
  sky130_fd_sc_hd__inv_2 _4595_ (
    .A(\g_bit[30].g_word[3].r_bit.Q ),
    .Y(_2233_)
  );
  sky130_fd_sc_hd__nor3_2 _4596_ (
    .A(_2233_),
    .B(_0280_),
    .C(_0082_),
    .Y(_2234_)
  );
  sky130_fd_sc_hd__and3_2 _4597_ (
    .A(\g_bit[30].g_word[24].r_bit.Q ),
    .B(_0077_),
    .C(_0078_),
    .X(_2235_)
  );
  sky130_fd_sc_hd__a2111o_2 _4598_ (
    .A1(\g_bit[30].g_word[29].r_bit.Q ),
    .A2(_0075_),
    .B1(_2232_),
    .C1(_2234_),
    .D1(_2235_),
    .X(_2236_)
  );
  sky130_fd_sc_hd__and3_2 _4599_ (
    .A(\g_bit[30].g_word[27].r_bit.Q ),
    .B(_0093_),
    .C(_0260_),
    .X(_2237_)
  );
  sky130_fd_sc_hd__a221o_2 _4600_ (
    .A1(\g_bit[30].g_word[6].r_bit.Q ),
    .A2(_0089_),
    .B1(_0091_),
    .B2(\g_bit[30].g_word[1].r_bit.Q ),
    .C1(_2237_),
    .X(_2238_)
  );
  sky130_fd_sc_hd__inv_2 _4601_ (
    .A(\g_bit[30].g_word[23].r_bit.Q ),
    .Y(_2239_)
  );
  sky130_fd_sc_hd__inv_2 _4602_ (
    .A(\g_bit[30].g_word[10].r_bit.Q ),
    .Y(_2240_)
  );
  sky130_fd_sc_hd__or3_2 _4603_ (
    .A(_2240_),
    .B(_0016_),
    .C(_0048_),
    .X(_2241_)
  );
  sky130_fd_sc_hd__inv_2 _4604_ (
    .A(\g_bit[30].g_word[9].r_bit.Q ),
    .Y(_2242_)
  );
  sky130_fd_sc_hd__or3_2 _4605_ (
    .A(_2242_),
    .B(_0103_),
    .C(_0041_),
    .X(_2243_)
  );
  sky130_fd_sc_hd__inv_2 _4606_ (
    .A(\g_bit[30].g_word[8].r_bit.Q ),
    .Y(_2244_)
  );
  sky130_fd_sc_hd__or3_2 _4607_ (
    .A(_2244_),
    .B(_0106_),
    .C(_0011_),
    .X(_2245_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4608_ (
    .A1(_2239_),
    .A2(_0100_),
    .B1(_2241_),
    .C1(_2243_),
    .D1(_2245_),
    .Y(_2246_)
  );
  sky130_fd_sc_hd__inv_2 _4609_ (
    .A(\g_bit[30].g_word[22].r_bit.Q ),
    .Y(_2247_)
  );
  sky130_fd_sc_hd__inv_2 _4610_ (
    .A(\g_bit[30].g_word[16].r_bit.Q ),
    .Y(_2248_)
  );
  sky130_fd_sc_hd__or3_2 _4611_ (
    .A(_2248_),
    .B(_0046_),
    .C(_0026_),
    .X(_2249_)
  );
  sky130_fd_sc_hd__inv_2 _4612_ (
    .A(\g_bit[30].g_word[14].r_bit.Q ),
    .Y(_2250_)
  );
  sky130_fd_sc_hd__or3_2 _4613_ (
    .A(_2250_),
    .B(_0107_),
    .C(_0028_),
    .X(_2251_)
  );
  sky130_fd_sc_hd__inv_2 _4614_ (
    .A(\g_bit[30].g_word[18].r_bit.Q ),
    .Y(_2252_)
  );
  sky130_fd_sc_hd__or3_2 _4615_ (
    .A(_2252_),
    .B(_0118_),
    .C(_0018_),
    .X(_2253_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4616_ (
    .A1(_2247_),
    .A2(_0115_),
    .B1(_2249_),
    .C1(_2251_),
    .D1(_2253_),
    .Y(_2254_)
  );
  sky130_fd_sc_hd__or4_2 _4617_ (
    .A(_2236_),
    .B(_2238_),
    .C(_2246_),
    .D(_2254_),
    .X(_2255_)
  );
  sky130_fd_sc_hd__or4_2 _4618_ (
    .A(_2223_),
    .B(_2225_),
    .C(_2230_),
    .D(_2255_),
    .X(_2256_)
  );
  sky130_fd_sc_hd__buf_1 _4619_ (
    .A(_2256_),
    .X(\g_bit[30].r_rs1.D )
  );
  sky130_fd_sc_hd__a32o_2 _4620_ (
    .A1(\g_bit[30].g_word[30].r_bit.Q ),
    .A2(_0151_),
    .A3(_0153_),
    .B1(_0158_),
    .B2(\g_bit[30].g_word[28].r_bit.Q ),
    .X(_2257_)
  );
  sky130_fd_sc_hd__a221o_2 _4621_ (
    .A1(\g_bit[30].g_word[4].r_bit.Q ),
    .A2(_0142_),
    .B1(_0149_),
    .B2(\g_bit[30].g_word[26].r_bit.Q ),
    .C1(_2257_),
    .X(_2258_)
  );
  sky130_fd_sc_hd__a22o_2 _4622_ (
    .A1(\g_bit[30].g_word[5].r_bit.Q ),
    .A2(_0171_),
    .B1(_0178_),
    .B2(\g_bit[30].g_word[2].r_bit.Q ),
    .X(_2259_)
  );
  sky130_fd_sc_hd__a221o_2 _4623_ (
    .A1(\g_bit[30].g_word[25].r_bit.Q ),
    .A2(_0163_),
    .B1(_0167_),
    .B2(\g_bit[30].g_word[31].r_bit.Q ),
    .C1(_2259_),
    .X(_2260_)
  );
  sky130_fd_sc_hd__a22o_2 _4624_ (
    .A1(\g_bit[30].g_word[13].r_bit.Q ),
    .A2(_0182_),
    .B1(_0185_),
    .B2(\g_bit[30].g_word[15].r_bit.Q ),
    .X(_2261_)
  );
  sky130_fd_sc_hd__a22o_2 _4625_ (
    .A1(\g_bit[30].g_word[20].r_bit.Q ),
    .A2(_0188_),
    .B1(_0190_),
    .B2(\g_bit[30].g_word[11].r_bit.Q ),
    .X(_2262_)
  );
  sky130_fd_sc_hd__a22o_2 _4626_ (
    .A1(\g_bit[30].g_word[19].r_bit.Q ),
    .A2(_0193_),
    .B1(_0195_),
    .B2(\g_bit[30].g_word[21].r_bit.Q ),
    .X(_2263_)
  );
  sky130_fd_sc_hd__a22o_2 _4627_ (
    .A1(\g_bit[30].g_word[17].r_bit.Q ),
    .A2(_0198_),
    .B1(_0200_),
    .B2(\g_bit[30].g_word[12].r_bit.Q ),
    .X(_2264_)
  );
  sky130_fd_sc_hd__or4_2 _4628_ (
    .A(_2261_),
    .B(_2262_),
    .C(_2263_),
    .D(_2264_),
    .X(_2265_)
  );
  sky130_fd_sc_hd__nor3_2 _4629_ (
    .A(_2231_),
    .B(_0132_),
    .C(_0209_),
    .Y(_2266_)
  );
  sky130_fd_sc_hd__nor3_2 _4630_ (
    .A(_2233_),
    .B(_0309_),
    .C(_0294_),
    .Y(_2267_)
  );
  sky130_fd_sc_hd__and3_2 _4631_ (
    .A(\g_bit[30].g_word[24].r_bit.Q ),
    .B(_0206_),
    .C(_0207_),
    .X(_2268_)
  );
  sky130_fd_sc_hd__a2111o_2 _4632_ (
    .A1(\g_bit[30].g_word[29].r_bit.Q ),
    .A2(_0204_),
    .B1(_2266_),
    .C1(_2267_),
    .D1(_2268_),
    .X(_2269_)
  );
  sky130_fd_sc_hd__and3_2 _4633_ (
    .A(\g_bit[30].g_word[27].r_bit.Q ),
    .B(_0219_),
    .C(_0298_),
    .X(_2270_)
  );
  sky130_fd_sc_hd__a221o_2 _4634_ (
    .A1(\g_bit[30].g_word[6].r_bit.Q ),
    .A2(_0215_),
    .B1(_0217_),
    .B2(\g_bit[30].g_word[1].r_bit.Q ),
    .C1(_2270_),
    .X(_2271_)
  );
  sky130_fd_sc_hd__or3_2 _4635_ (
    .A(_2240_),
    .B(_0145_),
    .C(_0177_),
    .X(_2272_)
  );
  sky130_fd_sc_hd__or3_2 _4636_ (
    .A(_2242_),
    .B(_0227_),
    .C(_0170_),
    .X(_2273_)
  );
  sky130_fd_sc_hd__or3_2 _4637_ (
    .A(_2244_),
    .B(_0229_),
    .C(_0140_),
    .X(_2274_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4638_ (
    .A1(_2239_),
    .A2(_0225_),
    .B1(_2272_),
    .C1(_2273_),
    .D1(_2274_),
    .Y(_2275_)
  );
  sky130_fd_sc_hd__or3_2 _4639_ (
    .A(_2248_),
    .B(_0155_),
    .C(_0175_),
    .X(_2276_)
  );
  sky130_fd_sc_hd__or3_2 _4640_ (
    .A(_2250_),
    .B(_0230_),
    .C(_0157_),
    .X(_2277_)
  );
  sky130_fd_sc_hd__or3_2 _4641_ (
    .A(_2252_),
    .B(_0240_),
    .C(_0147_),
    .X(_2278_)
  );
  sky130_fd_sc_hd__o2111ai_2 _4642_ (
    .A1(_2247_),
    .A2(_0236_),
    .B1(_2276_),
    .C1(_2277_),
    .D1(_2278_),
    .Y(_2279_)
  );
  sky130_fd_sc_hd__or4_2 _4643_ (
    .A(_2269_),
    .B(_2271_),
    .C(_2275_),
    .D(_2279_),
    .X(_2280_)
  );
  sky130_fd_sc_hd__or4_2 _4644_ (
    .A(_2258_),
    .B(_2260_),
    .C(_2265_),
    .D(_2280_),
    .X(_2281_)
  );
  sky130_fd_sc_hd__buf_1 _4645_ (
    .A(_2281_),
    .X(\g_bit[30].r_rs2.D )
  );
  sky130_fd_sc_hd__or2b_2 _4646_ (
    .A(i_rd[2]),
    .B_N(i_rd[3]),
    .X(_2282_)
  );
  sky130_fd_sc_hd__buf_1 _4647_ (
    .A(_2282_),
    .X(_2283_)
  );
  sky130_fd_sc_hd__or3b_2 _4649_ (
    .A(w_wr_sel_rd4),
    .B(i_rd[1]),
    .C_N(i_rd[0]),
    .X(_2285_)
  );
  sky130_fd_sc_hd__or3b_2 _4651_ (
    .A(i_rd[0]),
    .B(w_wr_sel_rd4),
    .C_N(i_rd[1]),
    .X(_2286_)
  );
  sky130_fd_sc_hd__nand2_2 _4653_ (
    .A(i_rd[1]),
    .B(i_rd[0]),
    .Y(_2287_)
  );
  sky130_fd_sc_hd__or2_2 _4654_ (
    .A(w_wr_sel_rd4),
    .B(_2287_),
    .X(_2288_)
  );
  sky130_fd_sc_hd__nand2_2 _4656_ (
    .A(i_rd[2]),
    .B(i_rd[3]),
    .Y(_2289_)
  );
  sky130_fd_sc_hd__or2_2 _4660_ (
    .A(i_rd[2]),
    .B(i_rd[3]),
    .X(_2290_)
  );
  sky130_fd_sc_hd__buf_1 _4661_ (
    .A(_2290_),
    .X(_2291_)
  );
  sky130_fd_sc_hd__or3b_2 _4663_ (
    .A(w_wr_sel_nrd4),
    .B(i_rd[1]),
    .C_N(i_rd[0]),
    .X(_2293_)
  );
  sky130_fd_sc_hd__or3b_2 _4665_ (
    .A(i_rd[0]),
    .B(w_wr_sel_nrd4),
    .C_N(i_rd[1]),
    .X(_2294_)
  );
  sky130_fd_sc_hd__or2_2 _4667_ (
    .A(_2287_),
    .B(w_wr_sel_nrd4),
    .X(_2295_)
  );
  sky130_fd_sc_hd__buf_1 _4670_ (
    .A(_2296_),
    .X(_2297_)
  );















  sky130_fd_sc_hd__or2b_2 rd3_nor_rd2 (
    .A(i_rd[3]),
    .B_N(i_rd[2]),
    .X(_2296_)
  );
  sky130_fd_sc_hd__nand3_2 wr_sel_rd4 (
    .A(i_write),
    .B(i_reset_n),
    .C(i_rd[4]),
    .Y(w_wr_sel_rd4)
  );
  sky130_fd_sc_hd__nand3b_2 wr_sel_nrd4 (
    .A_N(i_rd[4]),
    .B(i_reset_n),
    .C(i_write),
    .Y(w_wr_sel_nrd4)
  );
  sky130_fd_sc_hd__or3_2 wr_sel_rd4_rd0_or_rd1 (
    .A(i_rd[1]),
    .B(i_rd[0]),
    .C(w_wr_sel_rd4),
    .X(w_wr_sel_rd4_rd0_or_rd1)
  );
  sky130_fd_sc_hd__or3_2 wr_sel_nrd4_rd0_or_rd1 (
    .A(i_rd[1]),
    .B(i_rd[0]),
    .C(w_wr_sel_nrd4),
    .X(w_wr_sel_nrd4_rd0_or_rd1)
  );
  sky130_fd_sc_hd__nor2_2 \word[1].DE (
    .A(_2291_),
    .B(_2293_),
    .Y(\g_bit[0].g_word[1].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[2].DE (
    .A(_2291_),
    .B(_2294_),
    .Y(\g_bit[0].g_word[2].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[3].DE (
    .A(_2291_),
    .B(_2295_),
    .Y(\g_bit[0].g_word[3].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[4].DE (
    .A(_2297_),
    .B(w_wr_sel_nrd4_rd0_or_rd1),
    .Y(\g_bit[0].g_word[4].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[5].DE (
    .A(_2293_),
    .B(_2297_),
    .Y(\g_bit[0].g_word[5].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[6].DE (
    .A(_2294_),
    .B(_2297_),
    .Y(\g_bit[0].g_word[6].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[7].DE (
    .A(_2295_),
    .B(_2297_),
    .Y(\g_bit[0].g_word[7].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[8].DE (
    .A(_2283_),
    .B(w_wr_sel_nrd4_rd0_or_rd1),
    .Y(\g_bit[0].g_word[8].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[9].DE (
    .A(_2283_),
    .B(_2293_),
    .Y(\g_bit[0].g_word[9].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[10].DE (
    .A(_2283_),
    .B(_2294_),
    .Y(\g_bit[0].g_word[10].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[11].DE (
    .A(_2283_),
    .B(_2295_),
    .Y(\g_bit[0].g_word[11].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[12].DE (
    .A(_2289_),
    .B(w_wr_sel_nrd4_rd0_or_rd1),
    .Y(\g_bit[0].g_word[12].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[13].DE (
    .A(_2289_),
    .B(_2293_),
    .Y(\g_bit[0].g_word[13].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[14].DE (
    .A(_2289_),
    .B(_2294_),
    .Y(\g_bit[0].g_word[14].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[15].DE (
    .A(_2289_),
    .B(_2295_),
    .Y(\g_bit[0].g_word[15].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[16].DE (
    .A(_2291_),
    .B(w_wr_sel_rd4_rd0_or_rd1),
    .Y(\g_bit[0].g_word[16].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[17].DE (
    .A(_2285_),
    .B(_2291_),
    .Y(\g_bit[0].g_word[17].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[18].DE (
    .A(_2286_),
    .B(_2291_),
    .Y(\g_bit[0].g_word[18].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[19].DE (
    .A(_2288_),
    .B(_2291_),
    .Y(\g_bit[0].g_word[19].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[20].DE (
    .A(_2297_),
    .B(w_wr_sel_rd4_rd0_or_rd1),
    .Y(\g_bit[0].g_word[20].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[21].DE (
    .A(_2285_),
    .B(_2297_),
    .Y(\g_bit[0].g_word[21].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[22].DE (
    .A(_2286_),
    .B(_2297_),
    .Y(\g_bit[0].g_word[22].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[23].DE (
    .A(_2288_),
    .B(_2297_),
    .Y(\g_bit[0].g_word[23].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[24].DE (
    .A(_2283_),
    .B(w_wr_sel_rd4_rd0_or_rd1),
    .Y(\g_bit[0].g_word[24].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[25].DE (
    .A(_2283_),
    .B(_2285_),
    .Y(\g_bit[0].g_word[25].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[26].DE (
    .A(_2283_),
    .B(_2286_),
    .Y(\g_bit[0].g_word[26].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[27].DE (
    .A(_2283_),
    .B(_2288_),
    .Y(\g_bit[0].g_word[27].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[28].DE (
    .A(_2289_),
    .B(w_wr_sel_rd4_rd0_or_rd1),
    .Y(\g_bit[0].g_word[28].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[29].DE (
    .A(_2285_),
    .B(_2289_),
    .Y(\g_bit[0].g_word[29].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[30].DE (
    .A(_2286_),
    .B(_2289_),
    .Y(\g_bit[0].g_word[30].r_bit.DE )
  );
  sky130_fd_sc_hd__nor2_2 \word[31].DE (
    .A(_2288_),
    .B(_2289_),
    .Y(\g_bit[0].g_word[31].r_bit.DE )
  );
  sky130_fd_sc_hd__buf_2 \obuf1[0] (
    .A(\g_bit[0].r_rs1.Q ),
    .X(o_data1[0])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[1] (
    .A(\g_bit[1].r_rs1.Q ),
    .X(o_data1[1])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[2] (
    .A(\g_bit[2].r_rs1.Q ),
    .X(o_data1[2])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[3] (
    .A(\g_bit[3].r_rs1.Q ),
    .X(o_data1[3])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[4] (
    .A(\g_bit[4].r_rs1.Q ),
    .X(o_data1[4])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[5] (
    .A(\g_bit[5].r_rs1.Q ),
    .X(o_data1[5])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[6] (
    .A(\g_bit[6].r_rs1.Q ),
    .X(o_data1[6])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[7] (
    .A(\g_bit[7].r_rs1.Q ),
    .X(o_data1[7])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[8] (
    .A(\g_bit[8].r_rs1.Q ),
    .X(o_data1[8])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[9] (
    .A(\g_bit[9].r_rs1.Q ),
    .X(o_data1[9])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[10] (
    .A(\g_bit[10].r_rs1.Q ),
    .X(o_data1[10])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[11] (
    .A(\g_bit[11].r_rs1.Q ),
    .X(o_data1[11])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[12] (
    .A(\g_bit[12].r_rs1.Q ),
    .X(o_data1[12])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[13] (
    .A(\g_bit[13].r_rs1.Q ),
    .X(o_data1[13])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[14] (
    .A(\g_bit[14].r_rs1.Q ),
    .X(o_data1[14])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[15] (
    .A(\g_bit[15].r_rs1.Q ),
    .X(o_data1[15])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[16] (
    .A(\g_bit[16].r_rs1.Q ),
    .X(o_data1[16])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[17] (
    .A(\g_bit[17].r_rs1.Q ),
    .X(o_data1[17])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[18] (
    .A(\g_bit[18].r_rs1.Q ),
    .X(o_data1[18])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[19] (
    .A(\g_bit[19].r_rs1.Q ),
    .X(o_data1[19])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[20] (
    .A(\g_bit[20].r_rs1.Q ),
    .X(o_data1[20])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[21] (
    .A(\g_bit[21].r_rs1.Q ),
    .X(o_data1[21])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[22] (
    .A(\g_bit[22].r_rs1.Q ),
    .X(o_data1[22])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[23] (
    .A(\g_bit[23].r_rs1.Q ),
    .X(o_data1[23])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[24] (
    .A(\g_bit[24].r_rs1.Q ),
    .X(o_data1[24])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[25] (
    .A(\g_bit[25].r_rs1.Q ),
    .X(o_data1[25])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[26] (
    .A(\g_bit[26].r_rs1.Q ),
    .X(o_data1[26])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[27] (
    .A(\g_bit[27].r_rs1.Q ),
    .X(o_data1[27])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[28] (
    .A(\g_bit[28].r_rs1.Q ),
    .X(o_data1[28])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[29] (
    .A(\g_bit[29].r_rs1.Q ),
    .X(o_data1[29])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[30] (
    .A(\g_bit[30].r_rs1.Q ),
    .X(o_data1[30])
  );
  sky130_fd_sc_hd__buf_2 \obuf1[31] (
    .A(\g_bit[31].r_rs1.Q ),
    .X(o_data1[31])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[0] (
    .A(\g_bit[0].r_rs2.Q ),
    .X(o_data2[0])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[1] (
    .A(\g_bit[1].r_rs2.Q ),
    .X(o_data2[1])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[2] (
    .A(\g_bit[2].r_rs2.Q ),
    .X(o_data2[2])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[3] (
    .A(\g_bit[3].r_rs2.Q ),
    .X(o_data2[3])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[4] (
    .A(\g_bit[4].r_rs2.Q ),
    .X(o_data2[4])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[5] (
    .A(\g_bit[5].r_rs2.Q ),
    .X(o_data2[5])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[6] (
    .A(\g_bit[6].r_rs2.Q ),
    .X(o_data2[6])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[7] (
    .A(\g_bit[7].r_rs2.Q ),
    .X(o_data2[7])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[8] (
    .A(\g_bit[8].r_rs2.Q ),
    .X(o_data2[8])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[9] (
    .A(\g_bit[9].r_rs2.Q ),
    .X(o_data2[9])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[10] (
    .A(\g_bit[10].r_rs2.Q ),
    .X(o_data2[10])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[11] (
    .A(\g_bit[11].r_rs2.Q ),
    .X(o_data2[11])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[12] (
    .A(\g_bit[12].r_rs2.Q ),
    .X(o_data2[12])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[13] (
    .A(\g_bit[13].r_rs2.Q ),
    .X(o_data2[13])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[14] (
    .A(\g_bit[14].r_rs2.Q ),
    .X(o_data2[14])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[15] (
    .A(\g_bit[15].r_rs2.Q ),
    .X(o_data2[15])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[16] (
    .A(\g_bit[16].r_rs2.Q ),
    .X(o_data2[16])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[17] (
    .A(\g_bit[17].r_rs2.Q ),
    .X(o_data2[17])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[18] (
    .A(\g_bit[18].r_rs2.Q ),
    .X(o_data2[18])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[19] (
    .A(\g_bit[19].r_rs2.Q ),
    .X(o_data2[19])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[20] (
    .A(\g_bit[20].r_rs2.Q ),
    .X(o_data2[20])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[21] (
    .A(\g_bit[21].r_rs2.Q ),
    .X(o_data2[21])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[22] (
    .A(\g_bit[22].r_rs2.Q ),
    .X(o_data2[22])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[23] (
    .A(\g_bit[23].r_rs2.Q ),
    .X(o_data2[23])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[24] (
    .A(\g_bit[24].r_rs2.Q ),
    .X(o_data2[24])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[25] (
    .A(\g_bit[25].r_rs2.Q ),
    .X(o_data2[25])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[26] (
    .A(\g_bit[26].r_rs2.Q ),
    .X(o_data2[26])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[27] (
    .A(\g_bit[27].r_rs2.Q ),
    .X(o_data2[27])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[28] (
    .A(\g_bit[28].r_rs2.Q ),
    .X(o_data2[28])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[29] (
    .A(\g_bit[29].r_rs2.Q ),
    .X(o_data2[29])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[30] (
    .A(\g_bit[30].r_rs2.Q ),
    .X(o_data2[30])
  );
  sky130_fd_sc_hd__buf_2 \obuf2[31] (
    .A(\g_bit[31].r_rs2.Q ),
    .X(o_data2[31])
  );
  sky130_fd_sc_hd__mux2_2 \rs1_mux[0] (
    .A0(\r_rs1[0].Q ),
    .A1(i_rs1[0]),
    .S(i_rs_valid),
    .X(rs1[0])
  );
  sky130_fd_sc_hd__mux2_2 \rs1_mux[1] (
    .A0(\r_rs1[1].Q ),
    .A1(i_rs1[1]),
    .S(i_rs_valid),
    .X(rs1[1])
  );
  sky130_fd_sc_hd__mux2_2 \rs1_mux[2] (
    .A0(\r_rs1[2].Q ),
    .A1(i_rs1[2]),
    .S(i_rs_valid),
    .X(rs1[2])
  );
  sky130_fd_sc_hd__mux2_2 \rs1_mux[3] (
    .A0(\r_rs1[3].Q ),
    .A1(i_rs1[3]),
    .S(i_rs_valid),
    .X(rs1[3])
  );
  sky130_fd_sc_hd__mux2_2 \rs1_mux[4] (
    .A0(\r_rs1[4].Q ),
    .A1(i_rs1[4]),
    .S(i_rs_valid),
    .X(rs1[4])
  );
  sky130_fd_sc_hd__mux2_2 \rs2_mux[0] (
    .A0(\r_rs2[0].Q ),
    .A1(i_rs2[0]),
    .S(i_rs_valid),
    .X(rs2[0])
  );
  sky130_fd_sc_hd__mux2_2 \rs2_mux[1] (
    .A0(\r_rs2[1].Q ),
    .A1(i_rs2[1]),
    .S(i_rs_valid),
    .X(rs2[1])
  );
  sky130_fd_sc_hd__mux2_2 \rs2_mux[2] (
    .A0(\r_rs2[2].Q ),
    .A1(i_rs2[2]),
    .S(i_rs_valid),
    .X(rs2[2])
  );
  sky130_fd_sc_hd__mux2_2 \rs2_mux[3] (
    .A0(\r_rs2[3].Q ),
    .A1(i_rs2[3]),
    .S(i_rs_valid),
    .X(rs2[3])
  );
  sky130_fd_sc_hd__mux2_2 \rs2_mux[4] (
    .A0(\r_rs2[4].Q ),
    .A1(i_rs2[4]),
    .S(i_rs_valid),
    .X(rs2[4])
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[0].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[0].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[0].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[0].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[0].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[0].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[0].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[0].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[0].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[0].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[0].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[0].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[0].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[0].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[0].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[0].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[0].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[0].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[0].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[0].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[0].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[0].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[0].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[0].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[0].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[0].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[0].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[0].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[0].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[0].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[0].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[0]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[0].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[0].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[0].r_rs1.D ),
    .Q(\g_bit[0].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[0].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[0].r_rs2.D ),
    .Q(\g_bit[0].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[10].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[10].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[10].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[10].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[10].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[10].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[10].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[10].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[10].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[10].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[10].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[10].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[10].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[10].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[10].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[10].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[10].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[10].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[10].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[10].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[10].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[10].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[10].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[10].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[10].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[10].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[10].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[10].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[10].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[10].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[10].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[10]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[10].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[10].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[10].r_rs1.D ),
    .Q(\g_bit[10].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[10].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[10].r_rs2.D ),
    .Q(\g_bit[10].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[11].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[11].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[11].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[11].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[11].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[11].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[11].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[11].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[11].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[11].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[11].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[11].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[11].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[11].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[11].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[11].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[11].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[11].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[11].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[11].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[11].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[11].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[11].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[11].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[11].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[11].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[11].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[11].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[11].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[11].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[11].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[11]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[11].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[11].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[11].r_rs1.D ),
    .Q(\g_bit[11].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[11].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[11].r_rs2.D ),
    .Q(\g_bit[11].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[12].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[12].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[12].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[12].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[12].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[12].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[12].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[12].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[12].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[12].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[12].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[12].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[12].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[12].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[12].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[12].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[12].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[12].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[12].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[12].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[12].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[12].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[12].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[12].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[12].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[12].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[12].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[12].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[12].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[12].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[12].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[12]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[12].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[12].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[12].r_rs1.D ),
    .Q(\g_bit[12].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[12].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[12].r_rs2.D ),
    .Q(\g_bit[12].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[13].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[13].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[13].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[13].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[13].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[13].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[13].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[13].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[13].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[13].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[13].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[13].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[13].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[13].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[13].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[13].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[13].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[13].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[13].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[13].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[13].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[13].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[13].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[13].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[13].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[13].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[13].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[13].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[13].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[13].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[13].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[13]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[13].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[13].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[13].r_rs1.D ),
    .Q(\g_bit[13].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[13].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[13].r_rs2.D ),
    .Q(\g_bit[13].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[14].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[14].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[14].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[14].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[14].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[14].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[14].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[14].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[14].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[14].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[14].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[14].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[14].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[14].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[14].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[14].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[14].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[14].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[14].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[14].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[14].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[14].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[14].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[14].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[14].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[14].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[14].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[14].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[14].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[14].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[14].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[14]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[14].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[14].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[14].r_rs1.D ),
    .Q(\g_bit[14].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[14].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[14].r_rs2.D ),
    .Q(\g_bit[14].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[15].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[15].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[15].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[15].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[15].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[15].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[15].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[15].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[15].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[15].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[15].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[15].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[15].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[15].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[15].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[15].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[15].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[15].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[15].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[15].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[15].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[15].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[15].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[15].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[15].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[15].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[15].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[15].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[15].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[15].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[15].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[15]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[15].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[15].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[15].r_rs1.D ),
    .Q(\g_bit[15].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[15].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[15].r_rs2.D ),
    .Q(\g_bit[15].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[16].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[16].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[16].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[16].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[16].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[16].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[16].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[16].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[16].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[16].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[16].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[16].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[16].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[16].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[16].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[16].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[16].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[16].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[16].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[16].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[16].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[16].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[16].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[16].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[16].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[16].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[16].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[16].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[16].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[16].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[16].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[16]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[16].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[16].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[16].r_rs1.D ),
    .Q(\g_bit[16].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[16].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[16].r_rs2.D ),
    .Q(\g_bit[16].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[17].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[17].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[17].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[17].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[17].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[17].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[17].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[17].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[17].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[17].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[17].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[17].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[17].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[17].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[17].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[17].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[17].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[17].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[17].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[17].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[17].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[17].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[17].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[17].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[17].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[17].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[17].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[17].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[17].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[17].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[17].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[17]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[17].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[17].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[17].r_rs1.D ),
    .Q(\g_bit[17].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[17].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[17].r_rs2.D ),
    .Q(\g_bit[17].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[18].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[18].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[18].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[18].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[18].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[18].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[18].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[18].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[18].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[18].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[18].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[18].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[18].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[18].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[18].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[18].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[18].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[18].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[18].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[18].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[18].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[18].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[18].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[18].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[18].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[18].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[18].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[18].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[18].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[18].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[18].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[18]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[18].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[18].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[18].r_rs1.D ),
    .Q(\g_bit[18].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[18].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[18].r_rs2.D ),
    .Q(\g_bit[18].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[19].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[19].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[19].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[19].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[19].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[19].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[19].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[19].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[19].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[19].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[19].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[19].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[19].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[19].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[19].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[19].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[19].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[19].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[19].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[19].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[19].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[19].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[19].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[19].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[19].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[19].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[19].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[19].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[19].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[19].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[19].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[19]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[19].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[19].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[19].r_rs1.D ),
    .Q(\g_bit[19].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[19].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[19].r_rs2.D ),
    .Q(\g_bit[19].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[1].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[1].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[1].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[1].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[1].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[1].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[1].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[1].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[1].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[1].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[1].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[1].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[1].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[1].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[1].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[1].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[1].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[1].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[1].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[1].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[1].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[1].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[1].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[1].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[1].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[1].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[1].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[1].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[1].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[1].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[1].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[1]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[1].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[1].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[1].r_rs1.D ),
    .Q(\g_bit[1].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[1].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[1].r_rs2.D ),
    .Q(\g_bit[1].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[20].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[20].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[20].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[20].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[20].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[20].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[20].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[20].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[20].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[20].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[20].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[20].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[20].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[20].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[20].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[20].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[20].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[20].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[20].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[20].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[20].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[20].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[20].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[20].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[20].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[20].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[20].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[20].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[20].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[20].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[20].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[20]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[20].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[20].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[20].r_rs1.D ),
    .Q(\g_bit[20].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[20].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[20].r_rs2.D ),
    .Q(\g_bit[20].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[21].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[21].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[21].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[21].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[21].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[21].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[21].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[21].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[21].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[21].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[21].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[21].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[21].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[21].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[21].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[21].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[21].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[21].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[21].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[21].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[21].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[21].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[21].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[21].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[21].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[21].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[21].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[21].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[21].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[21].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[21].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[21]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[21].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[21].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[21].r_rs1.D ),
    .Q(\g_bit[21].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[21].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[21].r_rs2.D ),
    .Q(\g_bit[21].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[22].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[22].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[22].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[22].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[22].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[22].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[22].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[22].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[22].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[22].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[22].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[22].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[22].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[22].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[22].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[22].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[22].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[22].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[22].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[22].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[22].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[22].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[22].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[22].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[22].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[22].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[22].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[22].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[22].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[22].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[22].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[22]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[22].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[22].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[22].r_rs1.D ),
    .Q(\g_bit[22].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[22].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[22].r_rs2.D ),
    .Q(\g_bit[22].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[23].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[23].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[23].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[23].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[23].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[23].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[23].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[23].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[23].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[23].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[23].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[23].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[23].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[23].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[23].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[23].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[23].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[23].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[23].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[23].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[23].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[23].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[23].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[23].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[23].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[23].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[23].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[23].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[23].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[23].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[23].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[23]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[23].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[23].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[23].r_rs1.D ),
    .Q(\g_bit[23].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[23].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[23].r_rs2.D ),
    .Q(\g_bit[23].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[24].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[24].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[24].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[24].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[24].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[24].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[24].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[24].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[24].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[24].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[24].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[24].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[24].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[24].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[24].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[24].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[24].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[24].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[24].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[24].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[24].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[24].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[24].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[24].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[24].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[24].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[24].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[24].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[24].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[24].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[24].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[24]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[24].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[24].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[24].r_rs1.D ),
    .Q(\g_bit[24].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[24].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[24].r_rs2.D ),
    .Q(\g_bit[24].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[25].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[25].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[25].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[25].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[25].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[25].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[25].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[25].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[25].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[25].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[25].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[25].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[25].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[25].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[25].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[25].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[25].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[25].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[25].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[25].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[25].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[25].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[25].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[25].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[25].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[25].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[25].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[25].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[25].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[25].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[25].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[25]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[25].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[25].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[25].r_rs1.D ),
    .Q(\g_bit[25].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[25].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[25].r_rs2.D ),
    .Q(\g_bit[25].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[26].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[26].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[26].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[26].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[26].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[26].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[26].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[26].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[26].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[26].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[26].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[26].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[26].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[26].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[26].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[26].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[26].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[26].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[26].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[26].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[26].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[26].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[26].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[26].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[26].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[26].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[26].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[26].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[26].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[26].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[26].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[26]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[26].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[26].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[26].r_rs1.D ),
    .Q(\g_bit[26].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[26].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[26].r_rs2.D ),
    .Q(\g_bit[26].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[27].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[27].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[27].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[27].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[27].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[27].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[27].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[27].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[27].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[27].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[27].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[27].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[27].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[27].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[27].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[27].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[27].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[27].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[27].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[27].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[27].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[27].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[27].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[27].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[27].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[27].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[27].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[27].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[27].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[27].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[27].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[27]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[27].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[27].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[27].r_rs1.D ),
    .Q(\g_bit[27].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[27].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[27].r_rs2.D ),
    .Q(\g_bit[27].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[28].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[28].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[28].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[28].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[28].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[28].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[28].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[28].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[28].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[28].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[28].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[28].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[28].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[28].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[28].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[28].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[28].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[28].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[28].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[28].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[28].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[28].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[28].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[28].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[28].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[28].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[28].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[28].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[28].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[28].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[28].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[28]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[28].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[28].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[28].r_rs1.D ),
    .Q(\g_bit[28].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[28].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[28].r_rs2.D ),
    .Q(\g_bit[28].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[29].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[29].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[29].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[29].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[29].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[29].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[29].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[29].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[29].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[29].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[29].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[29].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[29].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[29].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[29].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[29].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[29].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[29].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[29].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[29].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[29].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[29].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[29].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[29].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[29].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[29].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[29].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[29].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[29].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[29].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[29].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[29]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[29].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[29].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[29].r_rs1.D ),
    .Q(\g_bit[29].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[29].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[29].r_rs2.D ),
    .Q(\g_bit[29].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[2].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[2].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[2].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[2].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[2].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[2].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[2].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[2].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[2].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[2].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[2].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[2].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[2].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[2].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[2].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[2].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[2].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[2].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[2].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[2].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[2].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[2].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[2].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[2].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[2].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[2].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[2].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[2].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[2].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[2].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[2].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[2]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[2].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[2].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[2].r_rs1.D ),
    .Q(\g_bit[2].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[2].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[2].r_rs2.D ),
    .Q(\g_bit[2].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[30].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[30].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[30].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[30].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[30].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[30].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[30].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[30].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[30].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[30].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[30].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[30].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[30].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[30].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[30].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[30].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[30].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[30].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[30].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[30].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[30].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[30].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[30].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[30].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[30].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[30].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[30].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[30].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[30].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[30].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[30].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[30]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[30].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[30].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[30].r_rs1.D ),
    .Q(\g_bit[30].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[30].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[30].r_rs2.D ),
    .Q(\g_bit[30].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[31].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[31].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[31].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[31].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[31].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[31].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[31].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[31].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[31].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[31].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[31].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[31].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[31].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[31].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[31].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[31].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[31].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[31].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[31].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[31].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[31].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[31].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[31].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[31].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[31].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[31].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[31].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[31].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[31].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[31].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[31].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[31]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[31].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[31].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[31].r_rs1.D ),
    .Q(\g_bit[31].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[31].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[31].r_rs2.D ),
    .Q(\g_bit[31].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[3].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[3].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[3].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[3].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[3].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[3].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[3].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[3].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[3].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[3].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[3].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[3].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[3].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[3].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[3].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[3].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[3].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[3].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[3].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[3].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[3].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[3].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[3].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[3].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[3].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[3].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[3].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[3].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[3].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[3].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[3].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[3]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[3].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[3].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[3].r_rs1.D ),
    .Q(\g_bit[3].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[3].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[3].r_rs2.D ),
    .Q(\g_bit[3].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[4].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[4].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[4].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[4].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[4].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[4].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[4].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[4].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[4].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[4].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[4].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[4].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[4].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[4].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[4].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[4].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[4].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[4].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[4].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[4].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[4].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[4].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[4].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[4].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[4].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[4].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[4].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[4].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[4].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[4].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[4].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[4]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[4].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[4].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[4].r_rs1.D ),
    .Q(\g_bit[4].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[4].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[4].r_rs2.D ),
    .Q(\g_bit[4].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[5].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[5].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[5].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[5].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[5].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[5].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[5].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[5].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[5].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[5].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[5].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[5].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[5].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[5].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[5].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[5].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[5].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[5].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[5].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[5].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[5].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[5].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[5].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[5].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[5].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[5].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[5].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[5].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[5].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[5].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[5].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[5]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[5].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[5].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[5].r_rs1.D ),
    .Q(\g_bit[5].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[5].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[5].r_rs2.D ),
    .Q(\g_bit[5].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[6].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[6].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[6].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[6].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[6].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[6].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[6].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[6].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[6].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[6].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[6].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[6].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[6].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[6].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[6].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[6].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[6].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[6].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[6].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[6].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[6].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[6].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[6].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[6].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[6].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[6].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[6].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[6].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[6].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[6].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[6].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[6]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[6].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[6].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[6].r_rs1.D ),
    .Q(\g_bit[6].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[6].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[6].r_rs2.D ),
    .Q(\g_bit[6].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[7].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[7].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[7].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[7].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[7].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[7].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[7].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[7].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[7].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[7].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[7].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[7].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[7].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[7].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[7].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[7].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[7].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[7].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[7].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[7].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[7].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[7].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[7].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[7].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[7].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[7].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[7].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[7].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[7].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[7].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[7].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[7]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[7].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[7].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[7].r_rs1.D ),
    .Q(\g_bit[7].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[7].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[7].r_rs2.D ),
    .Q(\g_bit[7].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[8].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[8].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[8].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[8].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[8].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[8].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[8].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[8].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[8].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[8].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[8].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[8].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[8].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[8].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[8].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[8].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[8].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[8].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[8].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[8].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[8].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[8].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[8].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[8].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[8].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[8].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[8].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[8].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[8].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[8].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[8].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[8]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[8].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[8].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[8].r_rs1.D ),
    .Q(\g_bit[8].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[8].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[8].r_rs2.D ),
    .Q(\g_bit[8].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[10].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[10].r_bit.DE ),
    .Q(\g_bit[9].g_word[10].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[11].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[11].r_bit.DE ),
    .Q(\g_bit[9].g_word[11].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[12].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[12].r_bit.DE ),
    .Q(\g_bit[9].g_word[12].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[13].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[13].r_bit.DE ),
    .Q(\g_bit[9].g_word[13].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[14].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[14].r_bit.DE ),
    .Q(\g_bit[9].g_word[14].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[15].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[15].r_bit.DE ),
    .Q(\g_bit[9].g_word[15].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[16].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[16].r_bit.DE ),
    .Q(\g_bit[9].g_word[16].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[17].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[17].r_bit.DE ),
    .Q(\g_bit[9].g_word[17].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[18].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[18].r_bit.DE ),
    .Q(\g_bit[9].g_word[18].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[19].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[19].r_bit.DE ),
    .Q(\g_bit[9].g_word[19].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[1].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[1].r_bit.DE ),
    .Q(\g_bit[9].g_word[1].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[20].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[20].r_bit.DE ),
    .Q(\g_bit[9].g_word[20].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[21].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[21].r_bit.DE ),
    .Q(\g_bit[9].g_word[21].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[22].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[22].r_bit.DE ),
    .Q(\g_bit[9].g_word[22].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[23].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[23].r_bit.DE ),
    .Q(\g_bit[9].g_word[23].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[24].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[24].r_bit.DE ),
    .Q(\g_bit[9].g_word[24].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[25].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[25].r_bit.DE ),
    .Q(\g_bit[9].g_word[25].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[26].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[26].r_bit.DE ),
    .Q(\g_bit[9].g_word[26].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[27].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[27].r_bit.DE ),
    .Q(\g_bit[9].g_word[27].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[28].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[28].r_bit.DE ),
    .Q(\g_bit[9].g_word[28].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[29].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[29].r_bit.DE ),
    .Q(\g_bit[9].g_word[29].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[2].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[2].r_bit.DE ),
    .Q(\g_bit[9].g_word[2].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[30].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[30].r_bit.DE ),
    .Q(\g_bit[9].g_word[30].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[31].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[31].r_bit.DE ),
    .Q(\g_bit[9].g_word[31].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[3].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[3].r_bit.DE ),
    .Q(\g_bit[9].g_word[3].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[4].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[4].r_bit.DE ),
    .Q(\g_bit[9].g_word[4].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[5].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[5].r_bit.DE ),
    .Q(\g_bit[9].g_word[5].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[6].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[6].r_bit.DE ),
    .Q(\g_bit[9].g_word[6].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[7].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[7].r_bit.DE ),
    .Q(\g_bit[9].g_word[7].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[8].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[8].r_bit.DE ),
    .Q(\g_bit[9].g_word[8].r_bit.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \g_bit[9].g_word[9].r_bit.r_bit  (
    .CLK(i_clk),
    .D(i_data[9]),
    .DE(\g_bit[0].g_word[9].r_bit.DE ),
    .Q(\g_bit[9].g_word[9].r_bit.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[9].r_rs1.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[9].r_rs1.D ),
    .Q(\g_bit[9].r_rs1.Q )
  );
  sky130_fd_sc_hd__dfxtp_1 \g_bit[9].r_rs2.r_bit  (
    .CLK(i_clk),
    .D(\g_bit[9].r_rs2.D ),
    .Q(\g_bit[9].r_rs2.Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \r_rs1[0].r_bit  (
    .CLK(i_clk),
    .D(i_rs1[0]),
    .DE(i_rs_valid),
    .Q(\r_rs1[0].Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \r_rs1[1].r_bit  (
    .CLK(i_clk),
    .D(i_rs1[1]),
    .DE(i_rs_valid),
    .Q(\r_rs1[1].Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \r_rs1[2].r_bit  (
    .CLK(i_clk),
    .D(i_rs1[2]),
    .DE(i_rs_valid),
    .Q(\r_rs1[2].Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \r_rs1[3].r_bit  (
    .CLK(i_clk),
    .D(i_rs1[3]),
    .DE(i_rs_valid),
    .Q(\r_rs1[3].Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \r_rs1[4].r_bit  (
    .CLK(i_clk),
    .D(i_rs1[4]),
    .DE(i_rs_valid),
    .Q(\r_rs1[4].Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \r_rs2[0].r_bit  (
    .CLK(i_clk),
    .D(i_rs2[0]),
    .DE(i_rs_valid),
    .Q(\r_rs2[0].Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \r_rs2[1].r_bit  (
    .CLK(i_clk),
    .D(i_rs2[1]),
    .DE(i_rs_valid),
    .Q(\r_rs2[1].Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \r_rs2[2].r_bit  (
    .CLK(i_clk),
    .D(i_rs2[2]),
    .DE(i_rs_valid),
    .Q(\r_rs2[2].Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \r_rs2[3].r_bit  (
    .CLK(i_clk),
    .D(i_rs2[3]),
    .DE(i_rs_valid),
    .Q(\r_rs2[3].Q )
  );
  sky130_fd_sc_hd__edfxtp_1 \r_rs2[4].r_bit  (
    .CLK(i_clk),
    .D(i_rs2[4]),
    .DE(i_rs_valid),
    .Q(\r_rs2[4].Q )
  );
endmodule
